----------------------------------------------------------------------------------
--
-- File retrieved, on 07/02/2010, from :
-- http://sebastien-viardot.imag.fr/Enseignements/Archi1A2s/sources/ROMPROG.vhd
--
-- Slightly altered to get rid of vendor-specific packages and adjust formatting
-- Now auto-filled by asrom script
--
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROMPROG is
  Port ( AD : in  STD_LOGIC_VECTOR (12 downto 0);
         D : out  STD_LOGIC_VECTOR (15 downto 0);
         CLK : in STD_LOGIC);
end ROMPROG;

architecture Behavioral of ROMPROG is
  constant low_address: natural := 0;
  constant high_address: natural := 8192;
  subtype octet is std_logic_vector( 15 downto 0 );
  type zone_memoire is
    array (natural range low_address to high_address-1) of octet;
  constant m: zone_memoire:= (
    0=>x"FFF7",	-- 1111111111110111  liw	r7, IRQ_mask
    1=>x"2000",	-- 0010000000000000  
    2=>x"F8C0",	-- 1111100011000000  bai	-, os_init
    3=>x"0100",	-- 0000000100000000  
   16=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_ack
   17=>x"2002",	-- 0010000000000010  
   18=>x"D001",	-- 1101000000000001  lw	r1, r0
   19=>x"F54A",	-- 1111010101001010  bspl	r2, r1, 5
   20=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_error
   21=>x"0050",	-- 0000000001010000  
   22=>x"F4CA",	-- 1111010011001010  bspl	r2, r1, 3
   23=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_kbd
   24=>x"0060",	-- 0000000001100000  
   25=>x"F40A",	-- 1111010000001010  bspl	r2, r1, 0
   26=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_tmr
   27=>x"0040",	-- 0000000001000000  
   28=>x"D201",	-- 1101001000000001  sw	r1, r0
   29=>x"FFFE",	-- 1111111111111110  reti
   64=>x"263F",	-- 0010011000111111  not r7, r7
   65=>x"D7C0",	-- 1101011111000000  out	r7
   66=>x"E383",	-- 1110001110000011  ba	-, r6
   80=>x"25FF",	-- 0010010111111111  xor	r7, r7, r7
   81=>x"D7C0",	-- 1101011111000000  out	r7
   82=>x"E383",	-- 1110001110000011  ba	-, r6
   96=>x"FFF2",	-- 1111111111110010  liw	r2, PS2_rx
   97=>x"2004",	-- 0010000000000100  
   98=>x"D012",	-- 1101000000010010  lw	r2, r2
   99=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map + 8
  100=>x"1808",	-- 0001100000001000  
  101=>x"D01B",	-- 1101000000011011  lw	r3, r3
  102=>x"1EBF",	-- 0001111010111111  mixll	r7, r7, r2
  103=>x"C784",	-- 1100011110000100  li	r4, 0xF0
  104=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  105=>x"8B20",	-- 1000101100100000  brieq	r4, int_kbd.release
  106=>x"C704",	-- 1100011100000100  li	r4, 0xE0
  107=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  108=>x"88E0",	-- 1000100011100000  brieq	r4, int_kbd.extended
  109=>x"FFF5",	-- 1111111111110101  liw	r5, paper_keys - 1
  110=>x"16BF",	-- 0001011010111111  
  111=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  112=>x"80E0",	-- 1000000011100000  brieq	r4, $+3
  113=>x"FFF5",	-- 1111111111110101  liw	r5, paper_keys + 10 - 1
  114=>x"16C9",	-- 0001011011001001  
  115=>x"042D",	-- 0000010000101101  inc	r5, r5
  116=>x"D02C",	-- 1101000000101100  lw	r4, r5
  117=>x"8560",	-- 1000010101100000  brieq	r4, scan_code_mismatch
  118=>x"6E24",	-- 0110111000100100  shr	r4, r4, 7
  119=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  120=>x"BEE4",	-- 1011111011100100  brine	r4, scan_code_loop
  121=>x"D02A",	-- 1101000000101010  lw	r2, r5
  122=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  123=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  124=>x"741B",	-- 0111010000011011  shr	r3, r3, 10
  125=>x"C00D",	-- 1100000000001101  li	r5, 1
  126=>x"0612",	-- 0000011000010010  dec	r2, r2
  127=>x"3AAA",	-- 0011101010101010  rrl	r2, r5, r2
  128=>x"FFF5",	-- 1111111111110101  liw	r5, key_press_map
  129=>x"1800",	-- 0001100000000000  
  130=>x"08ED",	-- 0000100011101101  add	r5, r5, r3
  131=>x"D02B",	-- 1101000000101011  lw	r3, r5
  132=>x"80E4",	-- 1000000011100100  brine	r4, scan_code_release
  133=>x"229B",	-- 0010001010011011  or	r3, r3, r2
  134=>x"80C3",	-- 1000000011000011  bri	-, scan_code_notify
  135=>x"2612",	-- 0010011000010010  not	r2, r2
  136=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  137=>x"D22B",	-- 1101001000101011  sw	r3, r5
  138=>x"C003",	-- 1100000000000011  li	r3, 0
  139=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  140=>x"1808",	-- 0001100000001000  
  141=>x"D223",	-- 1101001000100011  sw	r3, r4
  142=>x"E383",	-- 1110001110000011  ba	-, r6
  143=>x"C014",	-- 1100000000010100  li	r4, 2
  144=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  145=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  146=>x"1808",	-- 0001100000001000  
  147=>x"D223",	-- 1101001000100011  sw	r3, r4
  148=>x"E383",	-- 1110001110000011  ba	-, r6
  149=>x"C00C",	-- 1100000000001100  li	r4, 1
  150=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  151=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  152=>x"1808",	-- 0001100000001000  
  153=>x"D223",	-- 1101001000100011  sw	r3, r4
  154=>x"E383",	-- 1110001110000011  ba	-, r6
  256=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_mask
  257=>x"2000",	-- 0010000000000000  
  258=>x"C0C9",	-- 1100000011001001  li	r1, 0x19
  259=>x"D201",	-- 1101001000000001  sw	r1, r0
  260=>x"0400",	-- 0000010000000000  inc	r0, r0
  261=>x"CFF9",	-- 1100111111111001  li	r1, -1
  262=>x"D201",	-- 1101001000000001  sw	r1, r0
  263=>x"C03A",	-- 1100000000111010  li	r2, 7
  264=>x"0880",	-- 0000100010000000  add	r0, r0, r2
  265=>x"C0EA",	-- 1100000011101010  li	r2, 0x1D
  266=>x"D202",	-- 1101001000000010  sw	r2, r0
  267=>x"0400",	-- 0000010000000000  inc	r0, r0
  268=>x"C07A",	-- 1100000001111010  li	r2, 15
  269=>x"D202",	-- 1101001000000010  sw	r2, r0
  270=>x"FFF0",	-- 1111111111110000  liw	r0, key_press_map
  271=>x"1800",	-- 0001100000000000  
  272=>x"C001",	-- 1100000000000001  li	r1, 0
  273=>x"C042",	-- 1100000001000010  li	r2, 8
  274=>x"D201",	-- 1101001000000001  sw	r1, r0
  275=>x"0400",	-- 0000010000000000  inc	r0, r0
  276=>x"0612",	-- 0000011000010010  dec	r2, r2
  277=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  278=>x"C0F3",	-- 1100000011110011  li	r3, 30
  279=>x"CFFA",	-- 1100111111111010  li	r2, -1
  280=>x"D21A",	-- 1101001000011010  sw	r2, r3
  281=>x"8083",	-- 1000000010000011  bri	-, PaperGameStart
  282=>x"8003",	-- 1000000000000011  bri	-, PaperMenuLoop
  283=>x"FFF0",	-- 1111111111110000  liw	r0, paper_dir
  284=>x"1730",	-- 0001011100110000  
  285=>x"C001",	-- 1100000000000001  li	r1, 0
  286=>x"D201",	-- 1101001000000001  sw	r1, r0
  287=>x"0400",	-- 0000010000000000  inc	r0, r0
  288=>x"C4C1",	-- 1100010011000001  li	r1, 152
  289=>x"D201",	-- 1101001000000001  sw	r1, r0
  290=>x"0400",	-- 0000010000000000  inc	r0, r0
  291=>x"C001",	-- 1100000000000001  li	r1, 0
  292=>x"D201",	-- 1101001000000001  sw	r1, r0
  293=>x"0400",	-- 0000010000000000  inc	r0, r0
  294=>x"C401",	-- 1100010000000001  li	r1, 128
  295=>x"D201",	-- 1101001000000001  sw	r1, r0
  296=>x"0400",	-- 0000010000000000  inc	r0, r0
  297=>x"C001",	-- 1100000000000001  li	r1, 0
  298=>x"D201",	-- 1101001000000001  sw	r1, r0
  299=>x"0400",	-- 0000010000000000  inc	r0, r0
  300=>x"C0A1",	-- 1100000010100001  li	r1, 20
  301=>x"D201",	-- 1101001000000001  sw	r1, r0
  302=>x"0400",	-- 0000010000000000  inc	r0, r0
  303=>x"C029",	-- 1100000000101001  li	r1, 5
  304=>x"D201",	-- 1101001000000001  sw	r1, r0
  305=>x"0400",	-- 0000010000000000  inc	r0, r0
  306=>x"C000",	-- 1100000000000000  li	r0, 0
  307=>x"CFF9",	-- 1100111111111001  li	r1, -1
  308=>x"C0A2",	-- 1100000010100010  li	r2, 20
  309=>x"D201",	-- 1101001000000001  sw	r1, r0
  310=>x"0400",	-- 0000010000000000  inc	r0, r0
  311=>x"0612",	-- 0000011000010010  dec	r2, r2
  312=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  313=>x"C001",	-- 1100000000000001  li	r1, 0
  314=>x"FFF2",	-- 1111111111110010  liw	r2, 18*20
  315=>x"0168",	-- 0000000101101000  
  316=>x"D201",	-- 1101001000000001  sw	r1, r0
  317=>x"0400",	-- 0000010000000000  inc	r0, r0
  318=>x"0612",	-- 0000011000010010  dec	r2, r2
  319=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  320=>x"CFF9",	-- 1100111111111001  li	r1, -1
  321=>x"C0A2",	-- 1100000010100010  li	r2, 20
  322=>x"D201",	-- 1101001000000001  sw	r1, r0
  323=>x"0400",	-- 0000010000000000  inc	r0, r0
  324=>x"0612",	-- 0000011000010010  dec	r2, r2
  325=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  326=>x"C020",	-- 1100000000100000  li	r0, 4
  327=>x"C029",	-- 1100000000101001  li	r1, 5
  328=>x"FFF2",	-- 1111111111110010  liw	r2, paper_title
  329=>x"1738",	-- 0001011100111000  
  330=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  331=>x"0218",	-- 0000001000011000  
  332=>x"C790",	-- 1100011110010000  li	r0, 242
  333=>x"C009",	-- 1100000000001001  li	r1, 1
  334=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud
  335=>x"1720",	-- 0001011100100000  
  336=>x"C043",	-- 1100000001000011  li	r3, 8
  337=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  338=>x"02A3",	-- 0000001010100011  
  339=>x"C118",	-- 1100000100011000  li	r0, 35
  340=>x"C009",	-- 1100000000001001  li	r1, 1
  341=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  342=>x"173E",	-- 0001011100111110  
  343=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  344=>x"0218",	-- 0000001000011000  
  345=>x"C790",	-- 1100011110010000  li	r0, 242
  346=>x"C051",	-- 1100000001010001  li	r1, 10
  347=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud + 4
  348=>x"1724",	-- 0001011100100100  
  349=>x"C043",	-- 1100000001000011  li	r3, 8
  350=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  351=>x"02A3",	-- 0000001010100011  
  352=>x"C118",	-- 1100000100011000  li	r0, 35
  353=>x"C051",	-- 1100000001010001  li	r1, 10
  354=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  355=>x"173E",	-- 0001011100111110  
  356=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  357=>x"0218",	-- 0000001000011000  
  358=>x"FFF0",	-- 1111111111110000  liw	r0, 20*20
  359=>x"0190",	-- 0000000110010000  
  360=>x"C001",	-- 1100000000000001  li	r1, 0
  361=>x"FFF2",	-- 1111111111110010  liw	r2, 220*20
  362=>x"1130",	-- 0001000100110000  
  363=>x"D201",	-- 1101001000000001  sw	r1, r0
  364=>x"0400",	-- 0000010000000000  inc	r0, r0
  365=>x"0612",	-- 0000011000010010  dec	r2, r2
  366=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  367=>x"FFF3",	-- 1111111111110011  liw	r3, paper_dir
  368=>x"1730",	-- 0001011100110000  
  369=>x"D01C",	-- 1101000000011100  lw	r4, r3
  370=>x"041B",	-- 0000010000011011  inc	r3, r3
  371=>x"D018",	-- 1101000000011000  lw	r0, r3
  372=>x"041B",	-- 0000010000011011  inc	r3, r3
  373=>x"FFF2",	-- 1111111111110010  liw	r2, paper_sprites
  374=>x"16D0",	-- 0001011011010000  
  375=>x"4624",	-- 0100011000100100  shl	r4, r4, 3
  376=>x"0912",	-- 0000100100010010  add	r2, r2, r4
  377=>x"C083",	-- 1100000010000011  li	r3, 16
  378=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_16
  379=>x"0253",	-- 0000001001010011  
  380=>x"FFF2",	-- 1111111111110010  liw	r2, paper_dir
  381=>x"1730",	-- 0001011100110000  
  382=>x"D010",	-- 1101000000010000  lw	r0, r2
  383=>x"0412",	-- 0000010000010010  inc	r2, r2
  384=>x"D011",	-- 1101000000010001  lw	r1, r2
  385=>x"0600",	-- 0000011000000000  dec	r0, r0
  386=>x"80C4",	-- 1000000011000100  brine	r0, $+3
  387=>x"0609",	-- 0000011000001001  dec	r1, r1
  388=>x"8103",	-- 1000000100000011  bri	-, $+4
  389=>x"0600",	-- 0000011000000000  dec	r0, r0
  390=>x"8084",	-- 1000000010000100  brine	r0, $+2
  391=>x"0409",	-- 0000010000001001  inc	r1, r1
  392=>x"D211",	-- 1101001000010001  sw	r1, r2
  393=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  394=>x"1800",	-- 0001100000000000  
  395=>x"D01B",	-- 1101000000011011  lw	r3, r3
  396=>x"9718",	-- 1001011100011000  brieq	r3, event_not_kbd
  397=>x"F7DC",	-- 1111011111011100  bspl	r4, r3, 15
  398=>x"84A0",	-- 1000010010100000  brieq	r4, PaperGameQuit
  399=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  400=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveUp
  401=>x"F49C",	-- 1111010010011100  bspl	r4, r3, 2
  402=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveDOWN
  403=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  404=>x"8160",	-- 1000000101100000  brieq	r4, PaperNoMoveLEFT
  405=>x"FFF2",	-- 1111111111110010  liw	r2, paper_dir
  406=>x"1730",	-- 0001011100110000  
  407=>x"C010",	-- 1100000000010000  li	r0, 2
  408=>x"D210",	-- 1101001000010000  sw	r0, r2
  409=>x"F4DC",	-- 1111010011011100  bspl	r4, r3, 3
  410=>x"8160",	-- 1000000101100000  brieq	r4, PaperNoMoveRIGHT
  411=>x"FFF2",	-- 1111111111110010  liw	r2, paper_dir
  412=>x"1730",	-- 0001011100110000  
  413=>x"C008",	-- 1100000000001000  li	r0, 1
  414=>x"D210",	-- 1101001000010000  sw	r0, r2
  415=>x"B743",	-- 1011011101000011  bri	-, PaperGameLoop
  416=>x"FFFF",	-- 1111111111111111  reset
  417=>x"C040",	-- 1100000001000000  li	r0, 8
  418=>x"C041",	-- 1100000001000001  li	r1, 8
  419=>x"063F",	-- 0000011000111111  dec	r7, r7
  420=>x"D239",	-- 1101001000111001  sw	r1, r7
  421=>x"063F",	-- 0000011000111111  dec	r7, r7
  422=>x"D238",	-- 1101001000111000  sw	r0, r7
  423=>x"FFF2",	-- 1111111111110010  liw	r2, font_map + 4 * 0x23
  424=>x"134C",	-- 0001001101001100  
  425=>x"C043",	-- 1100000001000011  li	r3, 8
  426=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  427=>x"02A3",	-- 0000001010100011  
  428=>x"D038",	-- 1101000000111000  lw	r0, r7
  429=>x"043F",	-- 0000010000111111  inc	r7, r7
  430=>x"D039",	-- 1101000000111001  lw	r1, r7
  431=>x"043F",	-- 0000010000111111  inc	r7, r7
  432=>x"C0A2",	-- 1100000010100010  li	r2, 20
  433=>x"C003",	-- 1100000000000011  li	r3, 0
  434=>x"061B",	-- 0000011000011011  dec	r3, r3
  435=>x"BFDC",	-- 1011111111011100  brine	r3, $-1
  436=>x"0612",	-- 0000011000010010  dec	r2, r2
  437=>x"BF14",	-- 1011111100010100  brine	r2, $-4
  438=>x"FFF2",	-- 1111111111110010  liw	r2, key_press_map
  439=>x"1800",	-- 0001100000000000  
  440=>x"D012",	-- 1101000000010010  lw	r2, r2
  441=>x"8BD0",	-- 1000101111010000  brieq	r2, event_not_kbd
  442=>x"063F",	-- 0000011000111111  dec	r7, r7
  443=>x"D23A",	-- 1101001000111010  sw	r2, r7
  444=>x"063F",	-- 0000011000111111  dec	r7, r7
  445=>x"D239",	-- 1101001000111001  sw	r1, r7
  446=>x"063F",	-- 0000011000111111  dec	r7, r7
  447=>x"D238",	-- 1101001000111000  sw	r0, r7
  448=>x"FFF2",	-- 1111111111110010  liw	r2, font_map
  449=>x"12C0",	-- 0001001011000000  
  450=>x"C043",	-- 1100000001000011  li	r3, 8
  451=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  452=>x"02A3",	-- 0000001010100011  
  453=>x"D038",	-- 1101000000111000  lw	r0, r7
  454=>x"043F",	-- 0000010000111111  inc	r7, r7
  455=>x"D039",	-- 1101000000111001  lw	r1, r7
  456=>x"043F",	-- 0000010000111111  inc	r7, r7
  457=>x"D03A",	-- 1101000000111010  lw	r2, r7
  458=>x"043F",	-- 0000010000111111  inc	r7, r7
  459=>x"F413",	-- 1111010000010011  bspl	r3, r2, 0
  460=>x"81D8",	-- 1000000111011000  brieq	r3, event_kbd_no_up
  461=>x"C043",	-- 1100000001000011  li	r3, 8
  462=>x"0ACB",	-- 0000101011001011  sub	r3, r1, r3
  463=>x"809C",	-- 1000000010011100  brine	r3, event_kbd_no_clip_up
  464=>x"C781",	-- 1100011110000001  li	r1, 240
  465=>x"C043",	-- 1100000001000011  li	r3, 8
  466=>x"0AC9",	-- 0000101011001001  sub	r1, r1, r3
  467=>x"F453",	-- 1111010001010011  bspl	r3, r2, 1
  468=>x"8118",	-- 1000000100011000  brieq	r3, event_kbd_no_left
  469=>x"8084",	-- 1000000010000100  brine	r0, event_kbd_no_clip_left
  470=>x"C9C0",	-- 1100100111000000  li	r0, 39*8
  471=>x"0600",	-- 0000011000000000  dec	r0, r0
  472=>x"F493",	-- 1111010010010011  bspl	r3, r2, 2
  473=>x"81D8",	-- 1000000111011000  brieq	r3, event_kbd_no_down
  474=>x"C743",	-- 1100011101000011  li	r3, 232
  475=>x"0ACB",	-- 0000101011001011  sub	r3, r1, r3
  476=>x"809D",	-- 1000000010011101  brilt	r3, event_kbd_no_clip_down
  477=>x"C001",	-- 1100000000000001  li	r1, 0
  478=>x"C043",	-- 1100000001000011  li	r3, 8
  479=>x"08C9",	-- 0000100011001001  add	r1, r1, r3
  480=>x"F4D3",	-- 1111010011010011  bspl	r3, r2, 3
  481=>x"8198",	-- 1000000110011000  brieq	r3, event_kbd_no_right
  482=>x"C9C3",	-- 1100100111000011  li	r3, 39*8
  483=>x"0AC3",	-- 0000101011000011  sub	r3, r0, r3
  484=>x"809D",	-- 1000000010011101  brilt	r3, event_kbd_no_clip_right
  485=>x"CFF8",	-- 1100111111111000  li	r0, -1
  486=>x"0400",	-- 0000010000000000  inc	r0, r0
  487=>x"AF03",	-- 1010111100000011  bri	-, redraw
  488=>x"B383",	-- 1011001110000011  bri	-, event_loop
  489=>x"C750",	-- 1100011101010000  li	r0, 234
  490=>x"C1C2",	-- 1100000111000010  li	r2, 56
  491=>x"FAC6",	-- 1111101011000110  bail	-, r6, div_16_16
  492=>x"0201",	-- 0000001000000001  
  493=>x"C448",	-- 1100010001001000  li	r0, 137
  494=>x"C472",	-- 1100010001110010  li	r2, 142
  495=>x"FAC6",	-- 1111101011000110  bail	-, r6, mult_16_16
  496=>x"01F5",	-- 0000000111110101  
  497=>x"C03A",	-- 1100000000111010  li r2, 7
  498=>x"FAC6",	-- 1111101011000110  bail	-, r6, fact_16
  499=>x"020C",	-- 0000001000001100  
  500=>x"FFFF",	-- 1111111111111111  reset
  501=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  502=>x"2524",	-- 0010010100100100  xor	r4, r4, r4
  503=>x"C085",	-- 1100000010000101  li	r5, 16
  504=>x"0849",	-- 0000100001001001  add	r1, r1, r1
  505=>x"0C00",	-- 0000110000000000  adc	r0, r0, r0
  506=>x"0EDB",	-- 0000111011011011  sbc	r3, r3, r3
  507=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  508=>x"08C9",	-- 0000100011001001  add	r1, r1, r3
  509=>x"0D00",	-- 0000110100000000  adc	r0, r0, r4
  510=>x"062D",	-- 0000011000101101  dec	r5, r5
  511=>x"BE6C",	-- 1011111001101100  brine	r5, mult_16_16.loop
  512=>x"E383",	-- 1110001110000011  ba	-, r6
  513=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  514=>x"C084",	-- 1100000010000100  li	r4, 16
  515=>x"0800",	-- 0000100000000000  add	r0, r0, r0
  516=>x"0C49",	-- 0000110001001001  adc	r1, r1, r1
  517=>x"0A8B",	-- 0000101010001011  sub	r3, r1, r2
  518=>x"80DD",	-- 1000000011011101  brilt	r3, div_16_16.skip
  519=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  520=>x"0400",	-- 0000010000000000  inc	r0, r0
  521=>x"0624",	-- 0000011000100100  dec	r4, r4
  522=>x"BE64",	-- 1011111001100100  brine	r4, div_16_16.loop
  523=>x"E383",	-- 1110001110000011  ba	-, r6
  524=>x"2400",	-- 0010010000000000  xor	r0, r0, r0
  525=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  526=>x"8250",	-- 1000001001010000  brieq	r2, fact_16.end
  527=>x"0409",	-- 0000010000001001  inc	r1, r1
  528=>x"1008",	-- 0001000000001000  mova	r0, r1
  529=>x"FAC6",	-- 1111101011000110  bail	-, r6, mult_16_16
  530=>x"01F5",	-- 0000000111110101  
  531=>x"8104",	-- 1000000100000100  brine	r0, fact_16.overflow
  532=>x"01F5",	-- 0000000111110101  
  533=>x"0612",	-- 0000011000010010  dec	r2, r2
  534=>x"BE94",	-- 1011111010010100  brine	r2, fact_16.loop
  535=>x"E383",	-- 1110001110000011  ba	-, r6
  536=>x"063F",	-- 0000011000111111  dec	r7, r7
  537=>x"D23E",	-- 1101001000111110  sw	r6, r7
  538=>x"D013",	-- 1101000000010011  lw	r3, r2
  539=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  540=>x"84D8",	-- 1000010011011000  brieq	r3, puts.end
  541=>x"063F",	-- 0000011000111111  dec	r7, r7
  542=>x"D23A",	-- 1101001000111010  sw	r2, r7
  543=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  544=>x"0232",	-- 0000001000110010  
  545=>x"D03A",	-- 1101000000111010  lw	r2, r7
  546=>x"043F",	-- 0000010000111111  inc	r7, r7
  547=>x"D013",	-- 1101000000010011  lw	r3, r2
  548=>x"4E1B",	-- 0100111000011011  shl	r3, r3, 7
  549=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  550=>x"8258",	-- 1000001001011000  brieq	r3, puts.end
  551=>x"063F",	-- 0000011000111111  dec	r7, r7
  552=>x"D23A",	-- 1101001000111010  sw	r2, r7
  553=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  554=>x"0232",	-- 0000001000110010  
  555=>x"D03A",	-- 1101000000111010  lw	r2, r7
  556=>x"043F",	-- 0000010000111111  inc	r7, r7
  557=>x"0412",	-- 0000010000010010  inc	r2, r2
  558=>x"BB03",	-- 1011101100000011  bri	-, puts.loop
  559=>x"D03E",	-- 1101000000111110  lw	r6, r7
  560=>x"043F",	-- 0000010000111111  inc	r7, r7
  561=>x"E383",	-- 1110001110000011  ba	-, r6
  562=>x"063F",	-- 0000011000111111  dec	r7, r7
  563=>x"D23E",	-- 1101001000111110  sw	r6, r7
  564=>x"063F",	-- 0000011000111111  dec	r7, r7
  565=>x"D238",	-- 1101001000111000  sw	r0, r7
  566=>x"063F",	-- 0000011000111111  dec	r7, r7
  567=>x"D239",	-- 1101001000111001  sw	r1, r7
  568=>x"FFF2",	-- 1111111111110010  liw	r2, font_map
  569=>x"12C0",	-- 0001001011000000  
  570=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  571=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  572=>x"C043",	-- 1100000001000011  li	r3, 8
  573=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  574=>x"027D",	-- 0000001001111101  
  575=>x"D039",	-- 1101000000111001  lw	r1, r7
  576=>x"043F",	-- 0000010000111111  inc	r7, r7
  577=>x"D038",	-- 1101000000111000  lw	r0, r7
  578=>x"043F",	-- 0000010000111111  inc	r7, r7
  579=>x"0400",	-- 0000010000000000  inc	r0, r0
  580=>x"D03E",	-- 1101000000111110  lw	r6, r7
  581=>x"043F",	-- 0000010000111111  inc	r7, r7
  582=>x"E383",	-- 1110001110000011  ba	-, r6
  583=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  584=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  585=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  586=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  587=>x"C0A0",	-- 1100000010100000  li	r0, 20
  588=>x"D011",	-- 1101000000010001  lw	r1, r2
  589=>x"D221",	-- 1101001000100001  sw	r1, r4
  590=>x"0412",	-- 0000010000010010  inc	r2, r2
  591=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  592=>x"061B",	-- 0000011000011011  dec	r3, r3
  593=>x"BEDC",	-- 1011111011011100  brine	r3, put_sprite_16_aligned.loop
  594=>x"E383",	-- 1110001110000011  ba	-, r6
  595=>x"C07D",	-- 1100000001111101  li	r5, 15
  596=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  597=>x"6600",	-- 0110011000000000  shr	r0, r0, 3
  598=>x"BC68",	-- 1011110001101000  brieq	r5, put_sprite_16_aligned
  599=>x"062D",	-- 0000011000101101  dec	r5, r5
  600=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  601=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  602=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  603=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  604=>x"063F",	-- 0000011000111111  dec	r7, r7
  605=>x"D23B",	-- 1101001000111011  sw	r3, r7
  606=>x"D011",	-- 1101000000010001  lw	r1, r2
  607=>x"CFF8",	-- 1100111111111000  li	r0, -1
  608=>x"3D40",	-- 0011110101000000  rsr	r0, r0, r5
  609=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  610=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  611=>x"D023",	-- 1101000000100011  lw	r3, r4
  612=>x"2600",	-- 0010011000000000  not	r0, r0
  613=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  614=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  615=>x"D221",	-- 1101001000100001  sw	r1, r4
  616=>x"0424",	-- 0000010000100100  inc	r4, r4
  617=>x"D011",	-- 1101000000010001  lw	r1, r2
  618=>x"262D",	-- 0010011000101101  not	r5, r5
  619=>x"CFF8",	-- 1100111111111000  li	r0, -1
  620=>x"3F40",	-- 0011111101000000  rsl	r0, r0, r5
  621=>x"3B49",	-- 0011101101001001  rrl	r1, r1, r5
  622=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  623=>x"262D",	-- 0010011000101101  not	r5, r5
  624=>x"D023",	-- 1101000000100011  lw	r3, r4
  625=>x"2600",	-- 0010011000000000  not	r0, r0
  626=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  627=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  628=>x"D221",	-- 1101001000100001  sw	r1, r4
  629=>x"0412",	-- 0000010000010010  inc	r2, r2
  630=>x"C098",	-- 1100000010011000  li	r0, 19
  631=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  632=>x"D03B",	-- 1101000000111011  lw	r3, r7
  633=>x"043F",	-- 0000010000111111  inc	r7, r7
  634=>x"061B",	-- 0000011000011011  dec	r3, r3
  635=>x"B85C",	-- 1011100001011100  brine	r3, put_sprite_16.loop
  636=>x"E383",	-- 1110001110000011  ba	-, r6
  637=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  638=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  639=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  640=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  641=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  642=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  643=>x"C0A5",	-- 1100000010100101  li	r5, 20
  644=>x"8404",	-- 1000010000000100  brine	r0, put_sprite_8_aligned.loop1
  645=>x"D010",	-- 1101000000010000  lw	r0, r2
  646=>x"D021",	-- 1101000000100001  lw	r1, r4
  647=>x"1A41",	-- 0001101001000001  mixhl	r1, r0, r1
  648=>x"D221",	-- 1101001000100001  sw	r1, r4
  649=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  650=>x"061B",	-- 0000011000011011  dec	r3, r3
  651=>x"E398",	-- 1110001110011000  baeq	r3, r6
  652=>x"D021",	-- 1101000000100001  lw	r1, r4
  653=>x"1E41",	-- 0001111001000001  mixll	r1, r0, r1
  654=>x"D221",	-- 1101001000100001  sw	r1, r4
  655=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  656=>x"0412",	-- 0000010000010010  inc	r2, r2
  657=>x"061B",	-- 0000011000011011  dec	r3, r3
  658=>x"E398",	-- 1110001110011000  baeq	r3, r6
  659=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop0
  660=>x"D010",	-- 1101000000010000  lw	r0, r2
  661=>x"D021",	-- 1101000000100001  lw	r1, r4
  662=>x"1809",	-- 0001100000001001  mixhh	r1, r1, r0
  663=>x"D221",	-- 1101001000100001  sw	r1, r4
  664=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  665=>x"061B",	-- 0000011000011011  dec	r3, r3
  666=>x"E398",	-- 1110001110011000  baeq	r3, r6
  667=>x"D021",	-- 1101000000100001  lw	r1, r4
  668=>x"1A09",	-- 0001101000001001  mixhl	r1, r1, r0
  669=>x"D221",	-- 1101001000100001  sw	r1, r4
  670=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  671=>x"0412",	-- 0000010000010010  inc	r2, r2
  672=>x"061B",	-- 0000011000011011  dec	r3, r3
  673=>x"E398",	-- 1110001110011000  baeq	r3, r6
  674=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop1
  675=>x"C03D",	-- 1100000000111101  li	r5, 7
  676=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  677=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  678=>x"B5E8",	-- 1011010111101000  brieq	r5, put_sprite_8_aligned
  679=>x"062D",	-- 0000011000101101  dec	r5, r5
  680=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  681=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  682=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  683=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  684=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  685=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  686=>x"8A04",	-- 1000101000000100  brine	r0, put_sprite_8.loop1
  687=>x"D010",	-- 1101000000010000  lw	r0, r2
  688=>x"063F",	-- 0000011000111111  dec	r7, r7
  689=>x"D23A",	-- 1101001000111010  sw	r2, r7
  690=>x"C802",	-- 1100100000000010  li	r2, 0x100
  691=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  692=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  693=>x"D021",	-- 1101000000100001  lw	r1, r4
  694=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  695=>x"2612",	-- 0010011000010010  not	r2, r2
  696=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  697=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  698=>x"D221",	-- 1101001000100001  sw	r1, r4
  699=>x"C0A1",	-- 1100000010100001  li	r1, 20
  700=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  701=>x"D03A",	-- 1101000000111010  lw	r2, r7
  702=>x"043F",	-- 0000010000111111  inc	r7, r7
  703=>x"061B",	-- 0000011000011011  dec	r3, r3
  704=>x"E398",	-- 1110001110011000  baeq	r3, r6
  705=>x"D010",	-- 1101000000010000  lw	r0, r2
  706=>x"063F",	-- 0000011000111111  dec	r7, r7
  707=>x"D23A",	-- 1101001000111010  sw	r2, r7
  708=>x"1E00",	-- 0001111000000000  mixll	r0, r0, r0
  709=>x"C802",	-- 1100100000000010  li	r2, 0x100
  710=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  711=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  712=>x"D021",	-- 1101000000100001  lw	r1, r4
  713=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  714=>x"2612",	-- 0010011000010010  not	r2, r2
  715=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  716=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  717=>x"D221",	-- 1101001000100001  sw	r1, r4
  718=>x"C0A1",	-- 1100000010100001  li	r1, 20
  719=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  720=>x"D03A",	-- 1101000000111010  lw	r2, r7
  721=>x"043F",	-- 0000010000111111  inc	r7, r7
  722=>x"0412",	-- 0000010000010010  inc	r2, r2
  723=>x"061B",	-- 0000011000011011  dec	r3, r3
  724=>x"E398",	-- 1110001110011000  baeq	r3, r6
  725=>x"B683",	-- 1011011010000011  bri	-, put_sprite_8.loop0
  726=>x"D010",	-- 1101000000010000  lw	r0, r2
  727=>x"063F",	-- 0000011000111111  dec	r7, r7
  728=>x"D23A",	-- 1101001000111010  sw	r2, r7
  729=>x"063F",	-- 0000011000111111  dec	r7, r7
  730=>x"D23B",	-- 1101001000111011  sw	r3, r7
  731=>x"C802",	-- 1100100000000010  li	r2, 0x100
  732=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  733=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  734=>x"2080",	-- 0010000010000000  and	r0, r0, r2
  735=>x"D021",	-- 1101000000100001  lw	r1, r4
  736=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
  737=>x"261B",	-- 0010011000011011  not	r3, r3
  738=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  739=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
  740=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  741=>x"D221",	-- 1101001000100001  sw	r1, r4
  742=>x"0424",	-- 0000010000100100  inc	r4, r4
  743=>x"D021",	-- 1101000000100001  lw	r1, r4
  744=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  745=>x"261B",	-- 0010011000011011  not	r3, r3
  746=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  747=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
  748=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  749=>x"D221",	-- 1101001000100001  sw	r1, r4
  750=>x"C099",	-- 1100000010011001  li	r1, 19
  751=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  752=>x"D03B",	-- 1101000000111011  lw	r3, r7
  753=>x"043F",	-- 0000010000111111  inc	r7, r7
  754=>x"D03A",	-- 1101000000111010  lw	r2, r7
  755=>x"043F",	-- 0000010000111111  inc	r7, r7
  756=>x"061B",	-- 0000011000011011  dec	r3, r3
  757=>x"E398",	-- 1110001110011000  baeq	r3, r6
  758=>x"D010",	-- 1101000000010000  lw	r0, r2
  759=>x"4E00",	-- 0100111000000000  shl	r0, r0, 7
  760=>x"063F",	-- 0000011000111111  dec	r7, r7
  761=>x"D23A",	-- 1101001000111010  sw	r2, r7
  762=>x"063F",	-- 0000011000111111  dec	r7, r7
  763=>x"D23B",	-- 1101001000111011  sw	r3, r7
  764=>x"C802",	-- 1100100000000010  li	r2, 0x100
  765=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  766=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  767=>x"2080",	-- 0010000010000000  and	r0, r0, r2
  768=>x"D021",	-- 1101000000100001  lw	r1, r4
  769=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
  770=>x"261B",	-- 0010011000011011  not	r3, r3
  771=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  772=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
  773=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  774=>x"D221",	-- 1101001000100001  sw	r1, r4
  775=>x"0424",	-- 0000010000100100  inc	r4, r4
  776=>x"D021",	-- 1101000000100001  lw	r1, r4
  777=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  778=>x"261B",	-- 0010011000011011  not	r3, r3
  779=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  780=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
  781=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  782=>x"D221",	-- 1101001000100001  sw	r1, r4
  783=>x"C099",	-- 1100000010011001  li	r1, 19
  784=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  785=>x"D03B",	-- 1101000000111011  lw	r3, r7
  786=>x"043F",	-- 0000010000111111  inc	r7, r7
  787=>x"D03A",	-- 1101000000111010  lw	r2, r7
  788=>x"043F",	-- 0000010000111111  inc	r7, r7
  789=>x"0412",	-- 0000010000010010  inc	r2, r2
  790=>x"061B",	-- 0000011000011011  dec	r3, r3
  791=>x"E398",	-- 1110001110011000  baeq	r3, r6
  792=>x"AF83",	-- 1010111110000011  bri	-, put_sprite_8.loop1
    others => x"0000"
    );
begin
  process(CLK)
  begin
    if (CLK'event AND CLK='1') then
      D <= m(to_integer(unsigned(AD)));
    end if;
  end process;
end Behavioral;
