----------------------------------------------------------------------------------
--
-- File retrieved, on 07/02/2010, from :
-- http://sebastien-viardot.imag.fr/Enseignements/Archi1A2s/sources/ROMPROG.vhd
--
-- Slightly altered to get rid of vendor-specific packages and adjust formatting
-- Now auto-filled by asrom script
--
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROMPROG is
  Port ( AD : in  STD_LOGIC_VECTOR (12 downto 0);
         D : out  STD_LOGIC_VECTOR (15 downto 0);
         CLK : in STD_LOGIC);
end ROMPROG;

architecture Behavioral of ROMPROG is
  constant low_address: natural := 0;
  constant high_address: natural := 8192;
  subtype octet is std_logic_vector( 15 downto 0 );
  type zone_memoire is
    array (natural range low_address to high_address-1) of octet;
  constant m: zone_memoire:= (
    0=>x"FFF7",	-- 1111111111110111  liw	r7, IRQ_mask
    1=>x"2000",	-- 0010000000000000  
    2=>x"F8C0",	-- 1111100011000000  bai	-, os_init
    3=>x"0100",	-- 0000000100000000  
   16=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_ack
   17=>x"2002",	-- 0010000000000010  
   18=>x"D001",	-- 1101000000000001  lw	r1, r0
   19=>x"F54A",	-- 1111010101001010  bspl	r2, r1, 5
   20=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_error
   21=>x"0050",	-- 0000000001010000  
   22=>x"F4CA",	-- 1111010011001010  bspl	r2, r1, 3
   23=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_kbd
   24=>x"0060",	-- 0000000001100000  
   25=>x"F40A",	-- 1111010000001010  bspl	r2, r1, 0
   26=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_tmr
   27=>x"0040",	-- 0000000001000000  
   28=>x"D201",	-- 1101001000000001  sw	r1, r0
   29=>x"FFFE",	-- 1111111111111110  reti
   64=>x"263F",	-- 0010011000111111  not r7, r7
   65=>x"D7C0",	-- 1101011111000000  out	r7
   66=>x"E383",	-- 1110001110000011  ba	-, r6
   80=>x"25FF",	-- 0010010111111111  xor	r7, r7, r7
   81=>x"D7C0",	-- 1101011111000000  out	r7
   82=>x"E383",	-- 1110001110000011  ba	-, r6
   96=>x"FFF2",	-- 1111111111110010  liw	r2, PS2_rx
   97=>x"2004",	-- 0010000000000100  
   98=>x"D012",	-- 1101000000010010  lw	r2, r2
   99=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map + 8
  100=>x"16C8",	-- 0001011011001000  
  101=>x"D01B",	-- 1101000000011011  lw	r3, r3
  102=>x"1EBF",	-- 0001111010111111  mixll	r7, r7, r2
  103=>x"C784",	-- 1100011110000100  li	r4, 0xF0
  104=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  105=>x"8B20",	-- 1000101100100000  brieq	r4, int_kbd.release
  106=>x"C704",	-- 1100011100000100  li	r4, 0xE0
  107=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  108=>x"88E0",	-- 1000100011100000  brieq	r4, int_kbd.extended
  109=>x"FFF5",	-- 1111111111110101  liw	r5, paper_keys - 1
  110=>x"16CF",	-- 0001011011001111  
  111=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  112=>x"80E0",	-- 1000000011100000  brieq	r4, $+3
  113=>x"FFF5",	-- 1111111111110101  liw	r5, paper_keys + 11 - 1
  114=>x"16DA",	-- 0001011011011010  
  115=>x"042D",	-- 0000010000101101  inc	r5, r5
  116=>x"D02C",	-- 1101000000101100  lw	r4, r5
  117=>x"8560",	-- 1000010101100000  brieq	r4, scan_code_mismatch
  118=>x"6E24",	-- 0110111000100100  shr	r4, r4, 7
  119=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  120=>x"BEE4",	-- 1011111011100100  brine	r4, scan_code_loop
  121=>x"D02A",	-- 1101000000101010  lw	r2, r5
  122=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  123=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  124=>x"741B",	-- 0111010000011011  shr	r3, r3, 10
  125=>x"C00D",	-- 1100000000001101  li	r5, 1
  126=>x"0612",	-- 0000011000010010  dec	r2, r2
  127=>x"3AAA",	-- 0011101010101010  rrl	r2, r5, r2
  128=>x"FFF5",	-- 1111111111110101  liw	r5, key_press_map
  129=>x"16C0",	-- 0001011011000000  
  130=>x"08ED",	-- 0000100011101101  add	r5, r5, r3
  131=>x"D02B",	-- 1101000000101011  lw	r3, r5
  132=>x"80E4",	-- 1000000011100100  brine	r4, scan_code_release
  133=>x"229B",	-- 0010001010011011  or	r3, r3, r2
  134=>x"80C3",	-- 1000000011000011  bri	-, scan_code_notify
  135=>x"2612",	-- 0010011000010010  not	r2, r2
  136=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  137=>x"D22B",	-- 1101001000101011  sw	r3, r5
  138=>x"C003",	-- 1100000000000011  li	r3, 0
  139=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  140=>x"16C8",	-- 0001011011001000  
  141=>x"D223",	-- 1101001000100011  sw	r3, r4
  142=>x"E383",	-- 1110001110000011  ba	-, r6
  143=>x"C014",	-- 1100000000010100  li	r4, 2
  144=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  145=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  146=>x"16C8",	-- 0001011011001000  
  147=>x"D223",	-- 1101001000100011  sw	r3, r4
  148=>x"E383",	-- 1110001110000011  ba	-, r6
  149=>x"C00C",	-- 1100000000001100  li	r4, 1
  150=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  151=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  152=>x"16C8",	-- 0001011011001000  
  153=>x"D223",	-- 1101001000100011  sw	r3, r4
  154=>x"E383",	-- 1110001110000011  ba	-, r6
  256=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_mask
  257=>x"2000",	-- 0010000000000000  
  258=>x"C0C9",	-- 1100000011001001  li	r1, 0x19
  259=>x"D201",	-- 1101001000000001  sw	r1, r0
  260=>x"0400",	-- 0000010000000000  inc	r0, r0
  261=>x"CFF9",	-- 1100111111111001  li	r1, -1
  262=>x"D201",	-- 1101001000000001  sw	r1, r0
  263=>x"C03A",	-- 1100000000111010  li	r2, 7
  264=>x"0880",	-- 0000100010000000  add	r0, r0, r2
  265=>x"C0EA",	-- 1100000011101010  li	r2, 0x1D
  266=>x"D202",	-- 1101001000000010  sw	r2, r0
  267=>x"0400",	-- 0000010000000000  inc	r0, r0
  268=>x"C07A",	-- 1100000001111010  li	r2, 15
  269=>x"D202",	-- 1101001000000010  sw	r2, r0
  270=>x"0400",	-- 0000010000000000  inc	r0, r0
  271=>x"C0DA",	-- 1100000011011010  li	r2, 0x1B
  272=>x"D202",	-- 1101001000000010  sw	r2, r0
  273=>x"0400",	-- 0000010000000000  inc	r0, r0
  274=>x"FFF2",	-- 1111111111110010  liw	r2, 817
  275=>x"0331",	-- 0000001100110001  
  276=>x"D202",	-- 1101001000000010  sw	r2, r0
  277=>x"FFF0",	-- 1111111111110000  liw	r0, key_press_map
  278=>x"16C0",	-- 0001011011000000  
  279=>x"C001",	-- 1100000000000001  li	r1, 0
  280=>x"C042",	-- 1100000001000010  li	r2, 8
  281=>x"D201",	-- 1101001000000001  sw	r1, r0
  282=>x"0400",	-- 0000010000000000  inc	r0, r0
  283=>x"0612",	-- 0000011000010010  dec	r2, r2
  284=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  285=>x"8083",	-- 1000000010000011  bri	-, PaperGameStart
  286=>x"8003",	-- 1000000000000011  bri	-, PaperMenuLoop
  287=>x"FFF0",	-- 1111111111110000  liw	r0, paper_dir
  288=>x"179C",	-- 0001011110011100  
  289=>x"C001",	-- 1100000000000001  li	r1, 0
  290=>x"D201",	-- 1101001000000001  sw	r1, r0
  291=>x"0400",	-- 0000010000000000  inc	r0, r0
  292=>x"FFF1",	-- 1111111111110001  liw	r1, 152 * 8
  293=>x"04C0",	-- 0000010011000000  
  294=>x"D201",	-- 1101001000000001  sw	r1, r0
  295=>x"0400",	-- 0000010000000000  inc	r0, r0
  296=>x"C001",	-- 1100000000000001  li	r1, 0
  297=>x"D201",	-- 1101001000000001  sw	r1, r0
  298=>x"0400",	-- 0000010000000000  inc	r0, r0
  299=>x"FFF1",	-- 1111111111110001  liw	r1, 128 * 8
  300=>x"0400",	-- 0000010000000000  
  301=>x"D201",	-- 1101001000000001  sw	r1, r0
  302=>x"0400",	-- 0000010000000000  inc	r0, r0
  303=>x"C001",	-- 1100000000000001  li	r1, 0
  304=>x"D201",	-- 1101001000000001  sw	r1, r0
  305=>x"0400",	-- 0000010000000000  inc	r0, r0
  306=>x"C069",	-- 1100000001101001  li	r1, 13
  307=>x"D201",	-- 1101001000000001  sw	r1, r0
  308=>x"0400",	-- 0000010000000000  inc	r0, r0
  309=>x"C011",	-- 1100000000010001  li	r1, 2
  310=>x"D201",	-- 1101001000000001  sw	r1, r0
  311=>x"0400",	-- 0000010000000000  inc	r0, r0
  312=>x"FFF0",	-- 1111111111110000  liw	r0, paper_tilemap
  313=>x"17B0",	-- 0001011110110000  
  314=>x"C001",	-- 1100000000000001  li	r1, 0
  315=>x"C0C2",	-- 1100000011000010  li	r2, 6*4
  316=>x"D201",	-- 1101001000000001  sw	r1, r0
  317=>x"0400",	-- 0000010000000000  inc	r0, r0
  318=>x"0612",	-- 0000011000010010  dec	r2, r2
  319=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  320=>x"C000",	-- 1100000000000000  li	r0, 0
  321=>x"CFF9",	-- 1100111111111001  li	r1, -1
  322=>x"C0A2",	-- 1100000010100010  li	r2, 20
  323=>x"D201",	-- 1101001000000001  sw	r1, r0
  324=>x"0400",	-- 0000010000000000  inc	r0, r0
  325=>x"0612",	-- 0000011000010010  dec	r2, r2
  326=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  327=>x"C001",	-- 1100000000000001  li	r1, 0
  328=>x"FFF2",	-- 1111111111110010  liw	r2, 18*20
  329=>x"0168",	-- 0000000101101000  
  330=>x"D201",	-- 1101001000000001  sw	r1, r0
  331=>x"0400",	-- 0000010000000000  inc	r0, r0
  332=>x"0612",	-- 0000011000010010  dec	r2, r2
  333=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  334=>x"CFF9",	-- 1100111111111001  li	r1, -1
  335=>x"C0A2",	-- 1100000010100010  li	r2, 20
  336=>x"D201",	-- 1101001000000001  sw	r1, r0
  337=>x"0400",	-- 0000010000000000  inc	r0, r0
  338=>x"0612",	-- 0000011000010010  dec	r2, r2
  339=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  340=>x"C020",	-- 1100000000100000  li	r0, 4
  341=>x"C029",	-- 1100000000101001  li	r1, 5
  342=>x"FFF2",	-- 1111111111110010  liw	r2, paper_title
  343=>x"17A4",	-- 0001011110100100  
  344=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  345=>x"0298",	-- 0000001010011000  
  346=>x"C778",	-- 1100011101111000  li	r0, 239
  347=>x"C009",	-- 1100000000001001  li	r1, 1
  348=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud
  349=>x"1780",	-- 0001011110000000  
  350=>x"C043",	-- 1100000001000011  li	r3, 8
  351=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  352=>x"03A0",	-- 0000001110100000  
  353=>x"C0F8",	-- 1100000011111000  li	r0, 31
  354=>x"C009",	-- 1100000000001001  li	r1, 1
  355=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  356=>x"17A0",	-- 0001011110100000  
  357=>x"D012",	-- 1101000000010010  lw	r2, r2
  358=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum
  359=>x"02C7",	-- 0000001011000111  
  360=>x"C120",	-- 1100000100100000  li	r0, 36
  361=>x"C009",	-- 1100000000001001  li	r1, 1
  362=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  363=>x"17AA",	-- 0001011110101010  
  364=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  365=>x"0298",	-- 0000001010011000  
  366=>x"C778",	-- 1100011101111000  li	r0, 239
  367=>x"C051",	-- 1100000001010001  li	r1, 10
  368=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud + 4
  369=>x"1784",	-- 0001011110000100  
  370=>x"C043",	-- 1100000001000011  li	r3, 8
  371=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  372=>x"03A0",	-- 0000001110100000  
  373=>x"C0F8",	-- 1100000011111000  li	r0, 31
  374=>x"C051",	-- 1100000001010001  li	r1, 10
  375=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed + 1
  376=>x"17A1",	-- 0001011110100001  
  377=>x"D012",	-- 1101000000010010  lw	r2, r2
  378=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum
  379=>x"02C7",	-- 0000001011000111  
  380=>x"C120",	-- 1100000100100000  li	r0, 36
  381=>x"C051",	-- 1100000001010001  li	r1, 10
  382=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  383=>x"17AA",	-- 0001011110101010  
  384=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  385=>x"0298",	-- 0000001010011000  
  386=>x"FFF0",	-- 1111111111110000  liw	r0, 20*20
  387=>x"0190",	-- 0000000110010000  
  388=>x"C001",	-- 1100000000000001  li	r1, 0
  389=>x"FFF2",	-- 1111111111110010  liw	r2, 220*20
  390=>x"1130",	-- 0001000100110000  
  391=>x"D201",	-- 1101001000000001  sw	r1, r0
  392=>x"0400",	-- 0000010000000000  inc	r0, r0
  393=>x"0612",	-- 0000011000010010  dec	r2, r2
  394=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  395=>x"FFF5",	-- 1111111111110101  liw	r5, paper_tilemap
  396=>x"17B0",	-- 0001011110110000  
  397=>x"D02C",	-- 1101000000101100  lw	r4, r5
  398=>x"042D",	-- 0000010000101101  inc	r5, r5
  399=>x"8960",	-- 1000100101100000  brieq	r4, PaperGameTileSkip
  400=>x"063F",	-- 0000011000111111  dec	r7, r7
  401=>x"D23D",	-- 1101001000111101  sw	r5, r7
  402=>x"FFF3",	-- 1111111111110011  liw	r3, paper_tilemap
  403=>x"17B0",	-- 0001011110110000  
  404=>x"0AEB",	-- 0000101011101011  sub	r3, r5, r3
  405=>x"6E20",	-- 0110111000100000  shr	r0, r4, 7
  406=>x"6219",	-- 0110001000011001  shr	r1, r3, 1
  407=>x"4809",	-- 0100100000001001  shl	r1, r1, 4
  408=>x"C19A",	-- 1100000110011010  li	r2, 51
  409=>x"0889",	-- 0000100010001001  add	r1, r1, r2
  410=>x"FFF2",	-- 1111111111110010  liw	r2, paper_pos + 1
  411=>x"179E",	-- 0001011110011110  
  412=>x"D012",	-- 1101000000010010  lw	r2, r2
  413=>x"6412",	-- 0110010000010010  shr	r2, r2, 2
  414=>x"C0FB",	-- 1100000011111011  li	r3, 31
  415=>x"20D2",	-- 0010000011010010  and	r2, r2, r3
  416=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  417=>x"4E24",	-- 0100111000100100  shl	r4, r4, 7
  418=>x"6E24",	-- 0110111000100100  shr	r4, r4, 7
  419=>x"C00B",	-- 1100000000001011  li	r3, 1
  420=>x"FB06",	-- 1111101100000110  bailne	r0, r6, put_tile
  421=>x"0268",	-- 0000001001101000  
  422=>x"81E0",	-- 1000000111100000  brieq	r4, PaperGameSegmentSkip
  424=>x"C013",	-- 1100000000010011  li	r3, 2
  425=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_tile
  426=>x"0268",	-- 0000001001101000  
  427=>x"0624",	-- 0000011000100100  dec	r4, r4
  428=>x"BF64",	-- 1011111101100100  brine	r4, PaperGameSegmentLoop
  429=>x"C003",	-- 1100000000000011  li	r3, 0
  430=>x"C144",	-- 1100000101000100  li	r4, 40
  431=>x"0B04",	-- 0000101100000100  sub	r4, r0, r4
  432=>x"FB66",	-- 1111101101100110  baillt	r4, r6, put_tile
  433=>x"0268",	-- 0000001001101000  
  434=>x"D03D",	-- 1101000000111101  lw	r5, r7
  435=>x"043F",	-- 0000010000111111  inc	r7, r7
  436=>x"FFF4",	-- 1111111111110100  liw r4, paper_tilemap + 24
  437=>x"17C8",	-- 0001011111001000  
  438=>x"0B2C",	-- 0000101100101100  sub	r4, r5, r4
  439=>x"B5A5",	-- 1011010110100101  brilt	r4, PaperGameTileLoop
  440=>x"FFF3",	-- 1111111111110011  liw	r3, paper_speed
  441=>x"17A0",	-- 0001011110100000  
  442=>x"D01B",	-- 1101000000011011  lw	r3, r3
  443=>x"CF04",	-- 1100111100000100  li	r4, 0x1E0
  444=>x"211C",	-- 0010000100011100  and	r4, r3, r4
  445=>x"FFF3",	-- 1111111111110011  liw	r3, paper_pos
  446=>x"179D",	-- 0001011110011101  
  447=>x"D018",	-- 1101000000011000  lw	r0, r3
  448=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  449=>x"FFF2",	-- 1111111111110010  liw	r2, paper_sprites
  450=>x"1720",	-- 0001011100100000  
  451=>x"0912",	-- 0000100100010010  add	r2, r2, r4
  452=>x"C161",	-- 1100000101100001  li	r1, 44
  453=>x"C083",	-- 1100000010000011  li	r3, 16
  454=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_16_masked
  455=>x"0338",	-- 0000001100111000  
  456=>x"8FEC",	-- 1000111111101100  brine	r5, PaperGameFail
  458=>x"C028",	-- 1100000000101000  li	r0, 5
  459=>x"C001",	-- 1100000000000001  li	r1, 0
  460=>x"8043",	-- 1000000001000011  bri	-, $+1
  461=>x"0609",	-- 0000011000001001  dec	r1, r1
  462=>x"BF8C",	-- 1011111110001100  brine	r1, $-2
  463=>x"0600",	-- 0000011000000000  dec	r0, r0
  464=>x"BEC4",	-- 1011111011000100  brine	r0, $-5
  465=>x"FFF2",	-- 1111111111110010  liw	r2, paper_pos
  466=>x"179D",	-- 0001011110011101  
  467=>x"FFF3",	-- 1111111111110011  liw	r3, paper_speed
  468=>x"17A0",	-- 0001011110100000  
  469=>x"D010",	-- 1101000000010000  lw	r0, r2
  470=>x"D019",	-- 1101000000011001  lw	r1, r3
  471=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  472=>x"8BC5",	-- 1000101111000101  brilt	r0, PaperGameFail
  473=>x"FFF4",	-- 1111111111110100  liw	r4, 304*8
  474=>x"0980",	-- 0000100110000000  
  475=>x"0B04",	-- 0000101100000100  sub	r4, r0, r4
  476=>x"8AE1",	-- 1000101011100001  brige	r4, PaperGameFail
  477=>x"D210",	-- 1101001000010000  sw	r0, r2
  478=>x"0412",	-- 0000010000010010  inc	r2, r2
  479=>x"041B",	-- 0000010000011011  inc	r3, r3
  480=>x"D010",	-- 1101000000010000  lw	r0, r2
  481=>x"D019",	-- 1101000000011001  lw	r1, r3
  482=>x"C7FC",	-- 1100011111111100  li	r4, 0xFF
  483=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  484=>x"2101",	-- 0010000100000001  and	r1, r0, r4
  485=>x"D211",	-- 1101001000010001  sw	r1, r2
  486=>x"2624",	-- 0010011000100100  not	r4, r4
  487=>x"2100",	-- 0010000100000000  and	r0, r0, r4
  488=>x"FB06",	-- 1111101100000110  bailne	r0, r6, PaperMapScroll
  489=>x"0215",	-- 0000001000010101  
  490=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  491=>x"16C0",	-- 0001011011000000  
  492=>x"D01B",	-- 1101000000011011  lw	r3, r3
  493=>x"F818",	-- 1111100000011000  baieq	r3, PaperGameRedrawContent
  494=>x"0182",	-- 0000000110000010  
  495=>x"F7DC",	-- 1111011111011100  bspl	r4, r3, 15
  496=>x"8924",	-- 1000100100100100  brine	r4, PaperGameQuit
  497=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  498=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveUp
  499=>x"F49C",	-- 1111010010011100  bspl	r4, r3, 2
  500=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveDOWN
  501=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  502=>x"81E0",	-- 1000000111100000  brieq	r4, PaperNoMoveLEFT
  503=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  504=>x"17A0",	-- 0001011110100000  
  505=>x"D010",	-- 1101000000010000  lw	r0, r2
  506=>x"C02C",	-- 1100000000101100  li	r4, 5
  507=>x"0B00",	-- 0000101100000000  sub	r0, r0, r4
  508=>x"D210",	-- 1101001000010000  sw	r0, r2
  509=>x"F4DC",	-- 1111010011011100  bspl	r4, r3, 3
  510=>x"81E0",	-- 1000000111100000  brieq	r4, PaperNoMoveRIGHT
  511=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  512=>x"17A0",	-- 0001011110100000  
  513=>x"D010",	-- 1101000000010000  lw	r0, r2
  514=>x"C02C",	-- 1100000000101100  li	r4, 5
  515=>x"0900",	-- 0000100100000000  add	r0, r0, r4
  516=>x"D210",	-- 1101001000010000  sw	r0, r2
  517=>x"F8C0",	-- 1111100011000000  bai	-, PaperGameRedraw
  518=>x"0140",	-- 0000000101000000  
  519=>x"C000",	-- 1100000000000000  li	r0, 0
  520=>x"FFF2",	-- 1111111111110010  liw	r2, 240*20
  521=>x"12C0",	-- 0001001011000000  
  522=>x"D001",	-- 1101000000000001  lw	r1, r0
  523=>x"2609",	-- 0010011000001001  not	r1, r1
  524=>x"D201",	-- 1101001000000001  sw	r1, r0
  525=>x"0400",	-- 0000010000000000  inc	r0, r0
  526=>x"0612",	-- 0000011000010010  dec	r2, r2
  527=>x"BED4",	-- 1011111011010100  brine	r2, $-5
  528=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  529=>x"16C0",	-- 0001011011000000  
  530=>x"D01A",	-- 1101000000011010  lw	r2, r3
  531=>x"BFD0",	-- 1011111111010000  brieq	r2, $-1
  532=>x"FFFF",	-- 1111111111111111  reset
  533=>x"FFF0",	-- 1111111111110000  liw	r0, paper_tilemap
  534=>x"17B0",	-- 0001011110110000  
  535=>x"C021",	-- 1100000000100001  li	r1, 4
  536=>x"0841",	-- 0000100001000001  add	r1, r0, r1
  537=>x"C0A2",	-- 1100000010100010  li	r2, 5*4
  538=>x"D00B",	-- 1101000000001011  lw	r3, r1
  539=>x"D203",	-- 1101001000000011  sw	r3, r0
  540=>x"0400",	-- 0000010000000000  inc	r0, r0
  541=>x"0409",	-- 0000010000001001  inc	r1, r1
  542=>x"0612",	-- 0000011000010010  dec	r2, r2
  543=>x"BED4",	-- 1011111011010100  brine	r2, PaperGameScrollLoop
  544=>x"063F",	-- 0000011000111111  dec	r7, r7
  545=>x"D23E",	-- 1101001000111110  sw	r6, r7
  546=>x"FAC6",	-- 1111101011000110  bail	-, r6, rand16
  547=>x"0256",	-- 0000001001010110  
  548=>x"C02A",	-- 1100000000101010  li	r2, 0x05
  549=>x"208B",	-- 0010000010001011  and	r3, r1, r2
  550=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  551=>x"208C",	-- 0010000010001100  and	r4, r1, r2
  552=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  553=>x"1F19",	-- 0001111100011001  mixll	r1, r3, r4
  554=>x"D201",	-- 1101001000000001  sw	r1, r0
  555=>x"0400",	-- 0000010000000000  inc	r0, r0
  556=>x"C03A",	-- 1100000000111010  li	r2, 0x07
  557=>x"091C",	-- 0000100100011100  add r4, r3, r4
  558=>x"208B",	-- 0010000010001011  and	r3, r1, r2
  559=>x"091C",	-- 0000100100011100  add r4, r3, r4
  560=>x"C01B",	-- 1100000000011011  li	r3, 3
  561=>x"08E4",	-- 0000100011100100  add	r4, r4, r3
  562=>x"6209",	-- 0110001000001001  shr	r1, r1, 1
  563=>x"208B",	-- 0010000010001011  and	r3, r1, r2
  564=>x"091B",	-- 0000100100011011  add r3, r3, r4
  565=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  566=>x"208C",	-- 0010000010001100  and	r4, r1, r2
  567=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  568=>x"1F19",	-- 0001111100011001  mixll	r1, r3, r4
  569=>x"D201",	-- 1101001000000001  sw	r1, r0
  570=>x"0400",	-- 0000010000000000  inc	r0, r0
  571=>x"C02A",	-- 1100000000101010  li	r2, 0x05
  572=>x"091C",	-- 0000100100011100  add r4, r3, r4
  573=>x"208B",	-- 0010000010001011  and	r3, r1, r2
  574=>x"091C",	-- 0000100100011100  add r4, r3, r4
  575=>x"C01B",	-- 1100000000011011  li	r3, 3
  576=>x"08E4",	-- 0000100011100100  add	r4, r4, r3
  577=>x"6209",	-- 0110001000001001  shr	r1, r1, 1
  578=>x"208B",	-- 0010000010001011  and	r3, r1, r2
  579=>x"091B",	-- 0000100100011011  add r3, r3, r4
  580=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  581=>x"208C",	-- 0010000010001100  and	r4, r1, r2
  582=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  583=>x"1F19",	-- 0001111100011001  mixll	r1, r3, r4
  584=>x"D201",	-- 1101001000000001  sw	r1, r0
  585=>x"0400",	-- 0000010000000000  inc	r0, r0
  586=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed + 1
  587=>x"17A1",	-- 0001011110100001  
  588=>x"D011",	-- 1101000000010001  lw	r1, r2
  589=>x"0409",	-- 0000010000001001  inc	r1, r1
  590=>x"D211",	-- 1101001000010001  sw	r1, r2
  591=>x"D03E",	-- 1101000000111110  lw	r6, r7
  592=>x"043F",	-- 0000010000111111  inc	r7, r7
  593=>x"E383",	-- 1110001110000011  ba	-, r6
  594=>x"FFF2",	-- 1111111111110010  liw	r2, rand_seed
  595=>x"16C8",	-- 0001011011001000  
  596=>x"D210",	-- 1101001000010000  sw	r0, r2
  597=>x"E383",	-- 1110001110000011  ba	-, r6
  598=>x"FFF2",	-- 1111111111110010  liw	r2, rand_seed
  599=>x"16C8",	-- 0001011011001000  
  600=>x"D013",	-- 1101000000010011  lw	r3, r2
  601=>x"C7EC",	-- 1100011111101100  li	r4, 253
  602=>x"1F19",	-- 0001111100011001  mixll	r1, r3, r4
  603=>x"18E4",	-- 0001100011100100  mixhh	r4, r4, r3
  604=>x"C002",	-- 1100000000000010  li	r2, 0
  605=>x"0AC9",	-- 0000101011001001  sub	r1, r1, r3
  606=>x"0EA4",	-- 0000111010100100  sbc	r4, r4, r2
  607=>x"0EC9",	-- 0000111011001001  sbc	r1, r1, r3
  608=>x"0EA4",	-- 0000111010100100  sbc	r4, r4, r2
  609=>x"1B13",	-- 0001101100010011  mixhl	r3, r2, r4
  610=>x"0EC9",	-- 0000111011001001  sbc	r1, r1, r3
  611=>x"0C89",	-- 0000110010001001  adc	r1, r1, r2
  612=>x"FFF2",	-- 1111111111110010  liw	r2, rand_seed
  613=>x"16C8",	-- 0001011011001000  
  614=>x"D211",	-- 1101001000010001  sw	r1, r2
  615=>x"E383",	-- 1110001110000011  ba	-, r6
  616=>x"063F",	-- 0000011000111111  dec	r7, r7
  617=>x"D238",	-- 1101001000111000  sw	r0, r7
  618=>x"063F",	-- 0000011000111111  dec	r7, r7
  619=>x"D239",	-- 1101001000111001  sw	r1, r7
  620=>x"063F",	-- 0000011000111111  dec	r7, r7
  621=>x"D23A",	-- 1101001000111010  sw	r2, r7
  622=>x"063F",	-- 0000011000111111  dec	r7, r7
  623=>x"D23B",	-- 1101001000111011  sw	r3, r7
  624=>x"063F",	-- 0000011000111111  dec	r7, r7
  625=>x"D23C",	-- 1101001000111100  sw	r4, r7
  626=>x"063F",	-- 0000011000111111  dec	r7, r7
  627=>x"D23D",	-- 1101001000111101  sw	r5, r7
  628=>x"063F",	-- 0000011000111111  dec	r7, r7
  629=>x"D23E",	-- 1101001000111110  sw	r6, r7
  630=>x"FFF2",	-- 1111111111110010  liw	r2, paper_tiles
  631=>x"1790",	-- 0001011110010000  
  632=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  633=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  634=>x"C043",	-- 1100000001000011  li	r3, 8
  635=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  636=>x"037A",	-- 0000001101111010  
  637=>x"D03E",	-- 1101000000111110  lw	r6, r7
  638=>x"043F",	-- 0000010000111111  inc	r7, r7
  639=>x"D03D",	-- 1101000000111101  lw	r5, r7
  640=>x"043F",	-- 0000010000111111  inc	r7, r7
  641=>x"D03C",	-- 1101000000111100  lw	r4, r7
  642=>x"043F",	-- 0000010000111111  inc	r7, r7
  643=>x"D03B",	-- 1101000000111011  lw	r3, r7
  644=>x"043F",	-- 0000010000111111  inc	r7, r7
  645=>x"D03A",	-- 1101000000111010  lw	r2, r7
  646=>x"043F",	-- 0000010000111111  inc	r7, r7
  647=>x"D039",	-- 1101000000111001  lw	r1, r7
  648=>x"043F",	-- 0000010000111111  inc	r7, r7
  649=>x"D038",	-- 1101000000111000  lw	r0, r7
  650=>x"043F",	-- 0000010000111111  inc	r7, r7
  651=>x"0400",	-- 0000010000000000  inc	r0, r0
  652=>x"E383",	-- 1110001110000011  ba	-, r6
  653=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  654=>x"C084",	-- 1100000010000100  li	r4, 16
  655=>x"0800",	-- 0000100000000000  add	r0, r0, r0
  656=>x"0C49",	-- 0000110001001001  adc	r1, r1, r1
  657=>x"0A8B",	-- 0000101010001011  sub	r3, r1, r2
  658=>x"80DD",	-- 1000000011011101  brilt	r3, div_16_16.skip
  659=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  660=>x"0400",	-- 0000010000000000  inc	r0, r0
  661=>x"0624",	-- 0000011000100100  dec	r4, r4
  662=>x"BE64",	-- 1011111001100100  brine	r4, div_16_16.loop
  663=>x"E383",	-- 1110001110000011  ba	-, r6
  664=>x"063F",	-- 0000011000111111  dec	r7, r7
  665=>x"D23E",	-- 1101001000111110  sw	r6, r7
  666=>x"D013",	-- 1101000000010011  lw	r3, r2
  667=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  668=>x"84D8",	-- 1000010011011000  brieq	r3, puts.end
  669=>x"063F",	-- 0000011000111111  dec	r7, r7
  670=>x"D23A",	-- 1101001000111010  sw	r2, r7
  671=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  672=>x"02B2",	-- 0000001010110010  
  673=>x"D03A",	-- 1101000000111010  lw	r2, r7
  674=>x"043F",	-- 0000010000111111  inc	r7, r7
  675=>x"D013",	-- 1101000000010011  lw	r3, r2
  676=>x"4E1B",	-- 0100111000011011  shl	r3, r3, 7
  677=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  678=>x"8258",	-- 1000001001011000  brieq	r3, puts.end
  679=>x"063F",	-- 0000011000111111  dec	r7, r7
  680=>x"D23A",	-- 1101001000111010  sw	r2, r7
  681=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  682=>x"02B2",	-- 0000001010110010  
  683=>x"D03A",	-- 1101000000111010  lw	r2, r7
  684=>x"043F",	-- 0000010000111111  inc	r7, r7
  685=>x"0412",	-- 0000010000010010  inc	r2, r2
  686=>x"BB03",	-- 1011101100000011  bri	-, puts.loop
  687=>x"D03E",	-- 1101000000111110  lw	r6, r7
  688=>x"043F",	-- 0000010000111111  inc	r7, r7
  689=>x"E383",	-- 1110001110000011  ba	-, r6
  690=>x"063F",	-- 0000011000111111  dec	r7, r7
  691=>x"D23E",	-- 1101001000111110  sw	r6, r7
  692=>x"063F",	-- 0000011000111111  dec	r7, r7
  693=>x"D238",	-- 1101001000111000  sw	r0, r7
  694=>x"063F",	-- 0000011000111111  dec	r7, r7
  695=>x"D239",	-- 1101001000111001  sw	r1, r7
  696=>x"FFF2",	-- 1111111111110010  liw	r2, font_map
  697=>x"12C0",	-- 0001001011000000  
  698=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  699=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  700=>x"C043",	-- 1100000001000011  li	r3, 8
  701=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  702=>x"037A",	-- 0000001101111010  
  703=>x"D039",	-- 1101000000111001  lw	r1, r7
  704=>x"043F",	-- 0000010000111111  inc	r7, r7
  705=>x"D038",	-- 1101000000111000  lw	r0, r7
  706=>x"043F",	-- 0000010000111111  inc	r7, r7
  707=>x"0400",	-- 0000010000000000  inc	r0, r0
  708=>x"D03E",	-- 1101000000111110  lw	r6, r7
  709=>x"043F",	-- 0000010000111111  inc	r7, r7
  710=>x"E383",	-- 1110001110000011  ba	-, r6
  711=>x"063F",	-- 0000011000111111  dec	r7, r7
  712=>x"D23E",	-- 1101001000111110  sw	r6, r7
  713=>x"FFF4",	-- 1111111111110100  liw	r4, 10000
  714=>x"2710",	-- 0010011100010000  
  715=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  716=>x"02DA",	-- 0000001011011010  
  717=>x"FFF4",	-- 1111111111110100  liw	r4, 1000
  718=>x"03E8",	-- 0000001111101000  
  719=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  720=>x"02DA",	-- 0000001011011010  
  721=>x"C324",	-- 1100001100100100  li	r4, 100
  722=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  723=>x"02DA",	-- 0000001011011010  
  724=>x"C054",	-- 1100000001010100  li	r4, 10
  725=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  726=>x"02DA",	-- 0000001011011010  
  727=>x"D03E",	-- 1101000000111110  lw	r6, r7
  728=>x"043F",	-- 0000010000111111  inc	r7, r7
  729=>x"C00C",	-- 1100000000001100  li	r4, 1
  730=>x"C17B",	-- 1100000101111011  li	r3, 0x2F
  731=>x"041B",	-- 0000010000011011  inc	r3, r3
  732=>x"0B12",	-- 0000101100010010  sub	r2, r2, r4
  733=>x"BF91",	-- 1011111110010001  brige	r2, printnum.loop
  734=>x"0912",	-- 0000100100010010  add	r2, r2, r4
  735=>x"063F",	-- 0000011000111111  dec	r7, r7
  736=>x"D23E",	-- 1101001000111110  sw	r6, r7
  737=>x"063F",	-- 0000011000111111  dec	r7, r7
  738=>x"D23A",	-- 1101001000111010  sw	r2, r7
  739=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  740=>x"02B2",	-- 0000001010110010  
  741=>x"D03A",	-- 1101000000111010  lw	r2, r7
  742=>x"043F",	-- 0000010000111111  inc	r7, r7
  743=>x"D03E",	-- 1101000000111110  lw	r6, r7
  744=>x"043F",	-- 0000010000111111  inc	r7, r7
  745=>x"E383",	-- 1110001110000011  ba	-, r6
  746=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  747=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  748=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  749=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  750=>x"C0A0",	-- 1100000010100000  li	r0, 20
  751=>x"0412",	-- 0000010000010010  inc	r2, r2
  752=>x"D011",	-- 1101000000010001  lw	r1, r2
  753=>x"E421",	-- 1110010000100001  exw	r1, r4
  754=>x"0412",	-- 0000010000010010  inc	r2, r2
  755=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  756=>x"061B",	-- 0000011000011011  dec	r3, r3
  757=>x"BE9C",	-- 1011111010011100  brine	r3, put_sprite_16_aligned.loop
  758=>x"C005",	-- 1100000000000101  li	r5, 0
  759=>x"E383",	-- 1110001110000011  ba	-, r6
  760=>x"C07D",	-- 1100000001111101  li	r5, 15
  761=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  762=>x"6600",	-- 0110011000000000  shr	r0, r0, 3
  763=>x"BBE8",	-- 1011101111101000  brieq	r5, put_sprite_16_aligned
  764=>x"062D",	-- 0000011000101101  dec	r5, r5
  765=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  766=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  767=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  768=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  769=>x"063F",	-- 0000011000111111  dec	r7, r7
  770=>x"D23B",	-- 1101001000111011  sw	r3, r7
  771=>x"0412",	-- 0000010000010010  inc	r2, r2
  772=>x"D011",	-- 1101000000010001  lw	r1, r2
  773=>x"CFF8",	-- 1100111111111000  li	r0, -1
  774=>x"3D40",	-- 0011110101000000  rsr	r0, r0, r5
  775=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  776=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  777=>x"D023",	-- 1101000000100011  lw	r3, r4
  778=>x"2600",	-- 0010011000000000  not	r0, r0
  779=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  780=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  781=>x"E421",	-- 1110010000100001  exw	r1, r4
  782=>x"0424",	-- 0000010000100100  inc	r4, r4
  783=>x"D011",	-- 1101000000010001  lw	r1, r2
  784=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  785=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  786=>x"D023",	-- 1101000000100011  lw	r3, r4
  787=>x"2600",	-- 0010011000000000  not	r0, r0
  788=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  789=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  790=>x"E421",	-- 1110010000100001  exw	r1, r4
  791=>x"0412",	-- 0000010000010010  inc	r2, r2
  792=>x"C098",	-- 1100000010011000  li	r0, 19
  793=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  794=>x"D03B",	-- 1101000000111011  lw	r3, r7
  795=>x"043F",	-- 0000010000111111  inc	r7, r7
  796=>x"061B",	-- 0000011000011011  dec	r3, r3
  797=>x"B91C",	-- 1011100100011100  brine	r3, put_sprite_16.loop
  798=>x"C005",	-- 1100000000000101  li	r5, 0
  799=>x"E383",	-- 1110001110000011  ba	-, r6
  800=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  801=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  802=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  803=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  804=>x"C005",	-- 1100000000000101  li	r5, 0
  805=>x"D020",	-- 1101000000100000  lw	r0, r4
  806=>x"D011",	-- 1101000000010001  lw	r1, r2
  807=>x"0412",	-- 0000010000010010  inc	r2, r2
  808=>x"2040",	-- 0010000001000000  and	r0, r0, r1
  809=>x"D011",	-- 1101000000010001  lw	r1, r2
  810=>x"2240",	-- 0010001001000000  or	r0, r0, r1
  811=>x"E420",	-- 1110010000100000  exw	r0, r4
  812=>x"0612",	-- 0000011000010010  dec	r2, r2
  813=>x"D011",	-- 1101000000010001  lw	r1, r2
  814=>x"2609",	-- 0010011000001001  not	r1, r1
  815=>x"0412",	-- 0000010000010010  inc	r2, r2
  816=>x"2040",	-- 0010000001000000  and	r0, r0, r1
  817=>x"222D",	-- 0010001000101101  or	r5, r5, r0
  818=>x"0412",	-- 0000010000010010  inc	r2, r2
  819=>x"C0A0",	-- 1100000010100000  li	r0, 20
  820=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  821=>x"061B",	-- 0000011000011011  dec	r3, r3
  822=>x"AE5C",	-- 1010111001011100  brine	r3, put_sprite_16_aligned.loop
  823=>x"E383",	-- 1110001110000011  ba	-, r6
  824=>x"C07D",	-- 1100000001111101  li	r5, 15
  825=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  826=>x"6600",	-- 0110011000000000  shr	r0, r0, 3
  827=>x"B968",	-- 1011100101101000  brieq	r5, put_sprite_16_masked_aligned
  828=>x"062D",	-- 0000011000101101  dec	r5, r5
  829=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  830=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  831=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  832=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  833=>x"063F",	-- 0000011000111111  dec	r7, r7
  834=>x"D23E",	-- 1101001000111110  sw	r6, r7
  835=>x"102E",	-- 0001000000101110  mova	r6, r5
  836=>x"C005",	-- 1100000000000101  li	r5, 0
  837=>x"063F",	-- 0000011000111111  dec	r7, r7
  838=>x"D23B",	-- 1101001000111011  sw	r3, r7
  839=>x"063F",	-- 0000011000111111  dec	r7, r7
  840=>x"D23D",	-- 1101001000111101  sw	r5, r7
  841=>x"D010",	-- 1101000000010000  lw	r0, r2
  842=>x"3980",	-- 0011100110000000  rrr	r0, r0, r6
  843=>x"0412",	-- 0000010000010010  inc	r2, r2
  844=>x"D011",	-- 1101000000010001  lw	r1, r2
  845=>x"3989",	-- 0011100110001001  rrr	r1, r1, r6
  846=>x"CFFD",	-- 1100111111111101  li	r5, -1
  847=>x"3DAD",	-- 0011110110101101  rsr	r5, r5, r6
  848=>x"2149",	-- 0010000101001001  and	r1, r1, r5
  849=>x"D023",	-- 1101000000100011  lw	r3, r4
  850=>x"262D",	-- 0010011000101101  not	r5, r5
  851=>x"222D",	-- 0010001000101101  or	r5, r5, r0
  852=>x"215B",	-- 0010000101011011  and	r3, r3, r5
  853=>x"225B",	-- 0010001001011011  or	r3, r3, r1
  854=>x"E423",	-- 1110010000100011  exw	r3, r4
  855=>x"262D",	-- 0010011000101101  not	r5, r5
  856=>x"215B",	-- 0010000101011011  and	r3, r3, r5
  857=>x"D03D",	-- 1101000000111101  lw	r5, r7
  858=>x"043F",	-- 0000010000111111  inc	r7, r7
  859=>x"22ED",	-- 0010001011101101  or	r5, r5, r3
  860=>x"0424",	-- 0000010000100100  inc	r4, r4
  861=>x"063F",	-- 0000011000111111  dec	r7, r7
  862=>x"D23D",	-- 1101001000111101  sw	r5, r7
  863=>x"D011",	-- 1101000000010001  lw	r1, r2
  864=>x"3989",	-- 0011100110001001  rrr	r1, r1, r6
  865=>x"CFFD",	-- 1100111111111101  li	r5, -1
  866=>x"3DAD",	-- 0011110110101101  rsr	r5, r5, r6
  867=>x"262D",	-- 0010011000101101  not	r5, r5
  868=>x"2149",	-- 0010000101001001  and	r1, r1, r5
  869=>x"D023",	-- 1101000000100011  lw	r3, r4
  870=>x"262D",	-- 0010011000101101  not	r5, r5
  871=>x"222D",	-- 0010001000101101  or	r5, r5, r0
  872=>x"215B",	-- 0010000101011011  and	r3, r3, r5
  873=>x"225B",	-- 0010001001011011  or	r3, r3, r1
  874=>x"E423",	-- 1110010000100011  exw	r3, r4
  875=>x"262D",	-- 0010011000101101  not	r5, r5
  876=>x"215B",	-- 0010000101011011  and	r3, r3, r5
  877=>x"D03D",	-- 1101000000111101  lw	r5, r7
  878=>x"043F",	-- 0000010000111111  inc	r7, r7
  879=>x"22ED",	-- 0010001011101101  or	r5, r5, r3
  880=>x"0412",	-- 0000010000010010  inc	r2, r2
  881=>x"C098",	-- 1100000010011000  li	r0, 19
  882=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  883=>x"D03B",	-- 1101000000111011  lw	r3, r7
  884=>x"043F",	-- 0000010000111111  inc	r7, r7
  885=>x"061B",	-- 0000011000011011  dec	r3, r3
  886=>x"B3DC",	-- 1011001111011100  brine	r3, put_sprite_16_masked.loop
  887=>x"D03E",	-- 1101000000111110  lw	r6, r7
  888=>x"043F",	-- 0000010000111111  inc	r7, r7
  889=>x"E383",	-- 1110001110000011  ba	-, r6
  890=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  891=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  892=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  893=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  894=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  895=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  896=>x"C0A5",	-- 1100000010100101  li	r5, 20
  897=>x"8404",	-- 1000010000000100  brine	r0, put_sprite_8_aligned.loop1
  898=>x"D010",	-- 1101000000010000  lw	r0, r2
  899=>x"D021",	-- 1101000000100001  lw	r1, r4
  900=>x"1A41",	-- 0001101001000001  mixhl	r1, r0, r1
  901=>x"D221",	-- 1101001000100001  sw	r1, r4
  902=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  903=>x"061B",	-- 0000011000011011  dec	r3, r3
  904=>x"E398",	-- 1110001110011000  baeq	r3, r6
  905=>x"D021",	-- 1101000000100001  lw	r1, r4
  906=>x"1E41",	-- 0001111001000001  mixll	r1, r0, r1
  907=>x"D221",	-- 1101001000100001  sw	r1, r4
  908=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  909=>x"0412",	-- 0000010000010010  inc	r2, r2
  910=>x"061B",	-- 0000011000011011  dec	r3, r3
  911=>x"E398",	-- 1110001110011000  baeq	r3, r6
  912=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop0
  913=>x"D010",	-- 1101000000010000  lw	r0, r2
  914=>x"D021",	-- 1101000000100001  lw	r1, r4
  915=>x"1809",	-- 0001100000001001  mixhh	r1, r1, r0
  916=>x"D221",	-- 1101001000100001  sw	r1, r4
  917=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  918=>x"061B",	-- 0000011000011011  dec	r3, r3
  919=>x"E398",	-- 1110001110011000  baeq	r3, r6
  920=>x"D021",	-- 1101000000100001  lw	r1, r4
  921=>x"1A09",	-- 0001101000001001  mixhl	r1, r1, r0
  922=>x"D221",	-- 1101001000100001  sw	r1, r4
  923=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  924=>x"0412",	-- 0000010000010010  inc	r2, r2
  925=>x"061B",	-- 0000011000011011  dec	r3, r3
  926=>x"E398",	-- 1110001110011000  baeq	r3, r6
  927=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop1
  928=>x"C03D",	-- 1100000000111101  li	r5, 7
  929=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  930=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  931=>x"B5E8",	-- 1011010111101000  brieq	r5, put_sprite_8_aligned
  932=>x"062D",	-- 0000011000101101  dec	r5, r5
  933=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  934=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  935=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  936=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  937=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  938=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  939=>x"8A04",	-- 1000101000000100  brine	r0, put_sprite_8.loop1
  940=>x"D010",	-- 1101000000010000  lw	r0, r2
  941=>x"063F",	-- 0000011000111111  dec	r7, r7
  942=>x"D23A",	-- 1101001000111010  sw	r2, r7
  943=>x"C802",	-- 1100100000000010  li	r2, 0x100
  944=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  945=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  946=>x"D021",	-- 1101000000100001  lw	r1, r4
  947=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  948=>x"2612",	-- 0010011000010010  not	r2, r2
  949=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  950=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  951=>x"D221",	-- 1101001000100001  sw	r1, r4
  952=>x"C0A1",	-- 1100000010100001  li	r1, 20
  953=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  954=>x"D03A",	-- 1101000000111010  lw	r2, r7
  955=>x"043F",	-- 0000010000111111  inc	r7, r7
  956=>x"061B",	-- 0000011000011011  dec	r3, r3
  957=>x"E398",	-- 1110001110011000  baeq	r3, r6
  958=>x"D010",	-- 1101000000010000  lw	r0, r2
  959=>x"063F",	-- 0000011000111111  dec	r7, r7
  960=>x"D23A",	-- 1101001000111010  sw	r2, r7
  961=>x"1E00",	-- 0001111000000000  mixll	r0, r0, r0
  962=>x"C802",	-- 1100100000000010  li	r2, 0x100
  963=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  964=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  965=>x"D021",	-- 1101000000100001  lw	r1, r4
  966=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  967=>x"2612",	-- 0010011000010010  not	r2, r2
  968=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  969=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  970=>x"D221",	-- 1101001000100001  sw	r1, r4
  971=>x"C0A1",	-- 1100000010100001  li	r1, 20
  972=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  973=>x"D03A",	-- 1101000000111010  lw	r2, r7
  974=>x"043F",	-- 0000010000111111  inc	r7, r7
  975=>x"0412",	-- 0000010000010010  inc	r2, r2
  976=>x"061B",	-- 0000011000011011  dec	r3, r3
  977=>x"E398",	-- 1110001110011000  baeq	r3, r6
  978=>x"B683",	-- 1011011010000011  bri	-, put_sprite_8.loop0
  979=>x"D010",	-- 1101000000010000  lw	r0, r2
  980=>x"063F",	-- 0000011000111111  dec	r7, r7
  981=>x"D23A",	-- 1101001000111010  sw	r2, r7
  982=>x"063F",	-- 0000011000111111  dec	r7, r7
  983=>x"D23B",	-- 1101001000111011  sw	r3, r7
  984=>x"C802",	-- 1100100000000010  li	r2, 0x100
  985=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  986=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  987=>x"2080",	-- 0010000010000000  and	r0, r0, r2
  988=>x"D021",	-- 1101000000100001  lw	r1, r4
  989=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
  990=>x"261B",	-- 0010011000011011  not	r3, r3
  991=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  992=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
  993=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  994=>x"D221",	-- 1101001000100001  sw	r1, r4
  995=>x"0424",	-- 0000010000100100  inc	r4, r4
  996=>x"D021",	-- 1101000000100001  lw	r1, r4
  997=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  998=>x"261B",	-- 0010011000011011  not	r3, r3
  999=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
 1000=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
 1001=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
 1002=>x"D221",	-- 1101001000100001  sw	r1, r4
 1003=>x"C099",	-- 1100000010011001  li	r1, 19
 1004=>x"0864",	-- 0000100001100100  add	r4, r4, r1
 1005=>x"D03B",	-- 1101000000111011  lw	r3, r7
 1006=>x"043F",	-- 0000010000111111  inc	r7, r7
 1007=>x"D03A",	-- 1101000000111010  lw	r2, r7
 1008=>x"043F",	-- 0000010000111111  inc	r7, r7
 1009=>x"061B",	-- 0000011000011011  dec	r3, r3
 1010=>x"E398",	-- 1110001110011000  baeq	r3, r6
 1011=>x"D010",	-- 1101000000010000  lw	r0, r2
 1012=>x"4E00",	-- 0100111000000000  shl	r0, r0, 7
 1013=>x"063F",	-- 0000011000111111  dec	r7, r7
 1014=>x"D23A",	-- 1101001000111010  sw	r2, r7
 1015=>x"063F",	-- 0000011000111111  dec	r7, r7
 1016=>x"D23B",	-- 1101001000111011  sw	r3, r7
 1017=>x"C802",	-- 1100100000000010  li	r2, 0x100
 1018=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
 1019=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
 1020=>x"2080",	-- 0010000010000000  and	r0, r0, r2
 1021=>x"D021",	-- 1101000000100001  lw	r1, r4
 1022=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
 1023=>x"261B",	-- 0010011000011011  not	r3, r3
 1024=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
 1025=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
 1026=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
 1027=>x"D221",	-- 1101001000100001  sw	r1, r4
 1028=>x"0424",	-- 0000010000100100  inc	r4, r4
 1029=>x"D021",	-- 1101000000100001  lw	r1, r4
 1030=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
 1031=>x"261B",	-- 0010011000011011  not	r3, r3
 1032=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
 1033=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
 1034=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
 1035=>x"D221",	-- 1101001000100001  sw	r1, r4
 1036=>x"C099",	-- 1100000010011001  li	r1, 19
 1037=>x"0864",	-- 0000100001100100  add	r4, r4, r1
 1038=>x"D03B",	-- 1101000000111011  lw	r3, r7
 1039=>x"043F",	-- 0000010000111111  inc	r7, r7
 1040=>x"D03A",	-- 1101000000111010  lw	r2, r7
 1041=>x"043F",	-- 0000010000111111  inc	r7, r7
 1042=>x"0412",	-- 0000010000010010  inc	r2, r2
 1043=>x"061B",	-- 0000011000011011  dec	r3, r3
 1044=>x"E398",	-- 1110001110011000  baeq	r3, r6
 1045=>x"AF83",	-- 1010111110000011  bri	-, put_sprite_8.loop1
    others => x"0000"
    );
begin
  process(CLK)
  begin
    if (CLK'event AND CLK='1') then
      D <= m(to_integer(unsigned(AD)));
    end if;
  end process;
end Behavioral;
