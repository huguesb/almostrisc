----------------------------------------------------------------------------------
--
-- File retrieved, on 07/02/2010, from :
-- http://sebastien-viardot.imag.fr/Enseignements/Archi1A2s/sources/RAMDoublePort.vhd
--
-- Slightly altered to get rid of vendor-specific packages and adjust formatting
-- Now auto-filled by asrom script
--
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity RAMDoublePort is
    Port ( AD1 : in  STD_LOGIC_VECTOR (12 downto 0);
           AD2 : in  STD_LOGIC_VECTOR (12 downto 0);
           DIN1 : in  STD_LOGIC_VECTOR (15 downto 0);
           DOUT1 : out  STD_LOGIC_VECTOR (15 downto 0);
           WE1 : in  STD_LOGIC;
           DOUT2 : out  STD_LOGIC_VECTOR (15 downto 0);
           OE1 : in  STD_LOGIC;
           CE1 : in  STD_LOGIC;
			  CLK : in STD_LOGIC);
end RAMDoublePort;

 -- memory map :
 --     0 -  4799 : VGA-mapped RAM (320*240 pix, 16 pix per word => 4800 words)
 --  4800 -  5823 : font map (8*8 : 4 words per character, 256 chars => 1024 words)
 --  5824 -  8191 : user data (2368 words)

architecture Behavioral of RAMDoublePort is
 constant low_address: natural := 0;
 constant high_address: natural := 8192;  
 subtype octet is std_logic_vector( 15 downto 0 );
 type zone_memoire is
         array (natural range low_address to high_address) of octet;
 signal memoire: zone_memoire := (
  4804 => x"0050",
  4806 => x"8870",
  4808 => x"0050",
  4810 => x"7088",
  4812 => x"50F8",
  4813 => x"F8F8",
  4814 => x"F870",
  4815 => x"2000",
  4816 => x"2070",
  4817 => x"F8F8",
  4818 => x"F870",
  4819 => x"2000",
  4820 => x"7070",
  4821 => x"20F8",
  4822 => x"F820",
  4823 => x"7000",
  4824 => x"2070",
  4825 => x"F8F8",
  4826 => x"7020",
  4827 => x"7000",
  4829 => x"7070",
  4830 => x"7000",
  4832 => x"F8F8",
  4833 => x"8888",
  4834 => x"88F8",
  4835 => x"F800",
  4837 => x"7050",
  4838 => x"7000",
  4840 => x"F8F8",
  4841 => x"88A8",
  4842 => x"88F8",
  4843 => x"F800",
  4844 => x"2070",
  4845 => x"A820",
  4846 => x"7088",
  4847 => x"7000",
  4848 => x"7088",
  4849 => x"7020",
  4850 => x"20F8",
  4851 => x"2000",
  4852 => x"3838",
  4853 => x"2020",
  4854 => x"60E0",
  4855 => x"6000",
  4856 => x"7878",
  4857 => x"4858",
  4858 => x"58C0",
  4859 => x"C000",
  4860 => x"00A8",
  4861 => x"5088",
  4862 => x"50A8",
  4864 => x"4060",
  4865 => x"7078",
  4866 => x"7060",
  4867 => x"4000",
  4868 => x"1030",
  4869 => x"70F0",
  4870 => x"7030",
  4871 => x"1000",
  4872 => x"2070",
  4873 => x"A820",
  4874 => x"A870",
  4875 => x"2000",
  4876 => x"5050",
  4877 => x"5050",
  4878 => x"0050",
  4879 => x"5000",
  4880 => x"78E8",
  4881 => x"E878",
  4882 => x"2828",
  4883 => x"2800",
  4884 => x"78C8",
  4885 => x"A050",
  4886 => x"2898",
  4887 => x"F000",
  4890 => x"F8F8",
  4891 => x"F800",
  4892 => x"2070",
  4893 => x"2020",
  4894 => x"7020",
  4895 => x"F800",
  4896 => x"2070",
  4897 => x"F820",
  4898 => x"2020",
  4899 => x"2000",
  4900 => x"2020",
  4901 => x"2020",
  4902 => x"F870",
  4903 => x"2000",
  4904 => x"0020",
  4905 => x"30F8",
  4906 => x"3020",
  4908 => x"0020",
  4909 => x"60F8",
  4910 => x"6020",
  4913 => x"4078",
  4917 => x"50F8",
  4918 => x"5000",
  4920 => x"0020",
  4921 => x"2070",
  4922 => x"70F8",
  4923 => x"F800",
  4924 => x"F8F8",
  4925 => x"7070",
  4926 => x"2020",
  4932 => x"2020",
  4933 => x"2020",
  4934 => x"0020",
  4935 => x"2000",
  4936 => x"5050",
  4937 => x"5000",
  4940 => x"5050",
  4941 => x"F850",
  4942 => x"F850",
  4943 => x"5000",
  4944 => x"2070",
  4945 => x"A070",
  4946 => x"2870",
  4947 => x"2000",
  4948 => x"C0C8",
  4949 => x"1020",
  4950 => x"4098",
  4951 => x"1800",
  4952 => x"40A0",
  4953 => x"A040",
  4954 => x"A890",
  4955 => x"6800",
  4956 => x"2020",
  4957 => x"4000",
  4960 => x"1020",
  4961 => x"4040",
  4962 => x"4020",
  4963 => x"1000",
  4964 => x"4020",
  4965 => x"1010",
  4966 => x"1020",
  4967 => x"4000",
  4968 => x"A870",
  4969 => x"A800",
  4972 => x"0020",
  4973 => x"20F8",
  4974 => x"2020",
  4978 => x"6020",
  4979 => x"4000",
  4981 => x"00F8",
  4986 => x"0060",
  4987 => x"6000",
  4988 => x"0008",
  4989 => x"1020",
  4990 => x"4080",
  4992 => x"7088",
  4993 => x"98A8",
  4994 => x"C888",
  4995 => x"7000",
  4996 => x"20E0",
  4997 => x"2020",
  4998 => x"2020",
  4999 => x"F800",
  5000 => x"7088",
  5001 => x"0830",
  5002 => x"4080",
  5003 => x"F800",
  5004 => x"7088",
  5005 => x"0830",
  5006 => x"0888",
  5007 => x"7000",
  5008 => x"8888",
  5009 => x"88F8",
  5010 => x"0808",
  5011 => x"0800",
  5012 => x"F880",
  5013 => x"F008",
  5014 => x"0888",
  5015 => x"7000",
  5016 => x"7080",
  5017 => x"80F0",
  5018 => x"8888",
  5019 => x"7000",
  5020 => x"F808",
  5021 => x"0810",
  5022 => x"2020",
  5023 => x"2000",
  5024 => x"7088",
  5025 => x"8870",
  5026 => x"8888",
  5027 => x"7000",
  5028 => x"7088",
  5029 => x"8878",
  5030 => x"0808",
  5031 => x"7000",
  5032 => x"0060",
  5033 => x"6000",
  5034 => x"6060",
  5036 => x"0060",
  5037 => x"6000",
  5038 => x"6020",
  5039 => x"4000",
  5040 => x"1020",
  5041 => x"4080",
  5042 => x"4020",
  5043 => x"1000",
  5045 => x"F800",
  5046 => x"F800",
  5048 => x"4020",
  5049 => x"1008",
  5050 => x"1020",
  5051 => x"4000",
  5052 => x"7088",
  5053 => x"0810",
  5054 => x"2000",
  5055 => x"2000",
  5056 => x"7088",
  5057 => x"98A8",
  5058 => x"9880",
  5059 => x"7000",
  5060 => x"2020",
  5061 => x"5070",
  5062 => x"5088",
  5063 => x"8800",
  5064 => x"F088",
  5065 => x"88F0",
  5066 => x"8888",
  5067 => x"F000",
  5068 => x"7088",
  5069 => x"8080",
  5070 => x"8088",
  5071 => x"7000",
  5072 => x"F088",
  5073 => x"8888",
  5074 => x"8888",
  5075 => x"F000",
  5076 => x"F880",
  5077 => x"80F0",
  5078 => x"8080",
  5079 => x"F800",
  5080 => x"F880",
  5081 => x"80F0",
  5082 => x"8080",
  5083 => x"8000",
  5084 => x"7088",
  5085 => x"80B8",
  5086 => x"8888",
  5087 => x"7000",
  5088 => x"8888",
  5089 => x"88F8",
  5090 => x"8888",
  5091 => x"8800",
  5092 => x"F820",
  5093 => x"2020",
  5094 => x"2020",
  5095 => x"F800",
  5096 => x"0808",
  5097 => x"0808",
  5098 => x"0888",
  5099 => x"7000",
  5100 => x"8890",
  5101 => x"A0C0",
  5102 => x"A090",
  5103 => x"8800",
  5104 => x"8080",
  5105 => x"8080",
  5106 => x"8080",
  5107 => x"F800",
  5108 => x"88D8",
  5109 => x"A888",
  5110 => x"8888",
  5111 => x"8800",
  5112 => x"88C8",
  5113 => x"A898",
  5114 => x"8888",
  5115 => x"8800",
  5116 => x"7088",
  5117 => x"8888",
  5118 => x"8888",
  5119 => x"7000",
  5120 => x"F088",
  5121 => x"88F0",
  5122 => x"8080",
  5123 => x"8000",
  5124 => x"7088",
  5125 => x"8888",
  5126 => x"A890",
  5127 => x"6800",
  5128 => x"F088",
  5129 => x"88F0",
  5130 => x"9088",
  5131 => x"8800",
  5132 => x"7088",
  5133 => x"8070",
  5134 => x"0888",
  5135 => x"7000",
  5136 => x"F820",
  5137 => x"2020",
  5138 => x"2020",
  5139 => x"2000",
  5140 => x"8888",
  5141 => x"8888",
  5142 => x"8888",
  5143 => x"7000",
  5144 => x"8888",
  5145 => x"8888",
  5146 => x"8850",
  5147 => x"2000",
  5148 => x"8888",
  5149 => x"8888",
  5150 => x"A8D8",
  5151 => x"8800",
  5152 => x"8888",
  5153 => x"5020",
  5154 => x"5088",
  5155 => x"8800",
  5156 => x"8888",
  5157 => x"8850",
  5158 => x"2020",
  5159 => x"2000",
  5160 => x"F808",
  5161 => x"1020",
  5162 => x"4080",
  5163 => x"F800",
  5164 => x"7040",
  5165 => x"4040",
  5166 => x"4040",
  5167 => x"7000",
  5168 => x"0080",
  5169 => x"4020",
  5170 => x"1008",
  5172 => x"7010",
  5173 => x"1010",
  5174 => x"1010",
  5175 => x"7000",
  5176 => x"2050",
  5177 => x"8800",
  5183 => x"F800",
  5184 => x"0010",
  5185 => x"2000",
  5189 => x"7008",
  5190 => x"7888",
  5191 => x"7800",
  5192 => x"8080",
  5193 => x"80F0",
  5194 => x"8888",
  5195 => x"F000",
  5197 => x"7088",
  5198 => x"8088",
  5199 => x"7000",
  5200 => x"0808",
  5201 => x"0878",
  5202 => x"8888",
  5203 => x"7800",
  5205 => x"7088",
  5206 => x"F880",
  5207 => x"7800",
  5208 => x"3048",
  5209 => x"40E0",
  5210 => x"4040",
  5211 => x"4000",
  5213 => x"7888",
  5214 => x"7808",
  5215 => x"F000",
  5216 => x"8080",
  5217 => x"80F0",
  5218 => x"8888",
  5219 => x"8800",
  5220 => x"0020",
  5221 => x"0060",
  5222 => x"2020",
  5223 => x"7000",
  5224 => x"0010",
  5225 => x"0010",
  5226 => x"1090",
  5227 => x"6000",
  5228 => x"8080",
  5229 => x"90A0",
  5230 => x"C0A0",
  5231 => x"9800",
  5232 => x"6020",
  5233 => x"2020",
  5234 => x"2020",
  5235 => x"7000",
  5237 => x"D0A8",
  5238 => x"A888",
  5239 => x"8800",
  5241 => x"B0C8",
  5242 => x"8888",
  5243 => x"8800",
  5245 => x"7088",
  5246 => x"8888",
  5247 => x"7000",
  5249 => x"F088",
  5250 => x"F080",
  5251 => x"8000",
  5253 => x"7888",
  5254 => x"7808",
  5255 => x"0800",
  5257 => x"B0C8",
  5258 => x"8080",
  5259 => x"8000",
  5261 => x"7880",
  5262 => x"7008",
  5263 => x"F000",
  5264 => x"4040",
  5265 => x"E040",
  5266 => x"4048",
  5267 => x"3000",
  5269 => x"8888",
  5270 => x"8898",
  5271 => x"6800",
  5273 => x"8888",
  5274 => x"8850",
  5275 => x"2000",
  5277 => x"8888",
  5278 => x"88A8",
  5279 => x"5000",
  5281 => x"8850",
  5282 => x"2050",
  5283 => x"8800",
  5285 => x"8850",
  5286 => x"2040",
  5287 => x"8000",
  5289 => x"F810",
  5290 => x"2040",
  5291 => x"F800",
  5292 => x"1820",
  5293 => x"2040",
  5294 => x"2020",
  5295 => x"1800",
  5296 => x"2020",
  5297 => x"2000",
  5298 => x"2020",
  5299 => x"2000",
  5300 => x"6010",
  5301 => x"1008",
  5302 => x"1010",
  5303 => x"6000",
  5305 => x"40A8",
  5306 => x"1000",
  5308 => x"0020",
  5309 => x"5088",
  5310 => x"8888",
  5311 => x"F800",
  5312 => x"7088",
  5313 => x"8088",
  5314 => x"7020",
  5315 => x"C000",
  5316 => x"0070",
  5317 => x"8088",
  5318 => x"7020",
  5319 => x"C000",
  5320 => x"1448",
  5321 => x"88C8",
  5322 => x"A898",
  5323 => x"8800",
  5324 => x"2850",
  5325 => x"00B0",
  5326 => x"C888",
  5327 => x"8800",
  5328 => x"1020",
  5329 => x"7088",
  5330 => x"F888",
  5331 => x"8800",
  5332 => x"4020",
  5333 => x"7088",
  5334 => x"F888",
  5335 => x"8800",
  5336 => x"5000",
  5337 => x"7088",
  5338 => x"F888",
  5339 => x"8800",
  5340 => x"2050",
  5341 => x"0070",
  5342 => x"88F8",
  5343 => x"8800",
  5344 => x"1020",
  5345 => x"F880",
  5346 => x"F080",
  5347 => x"F800",
  5348 => x"4020",
  5349 => x"F880",
  5350 => x"F080",
  5351 => x"F800",
  5352 => x"5000",
  5353 => x"F880",
  5354 => x"F080",
  5355 => x"F800",
  5356 => x"2050",
  5357 => x"F880",
  5358 => x"F080",
  5359 => x"F800",
  5360 => x"1020",
  5361 => x"F820",
  5362 => x"2020",
  5363 => x"F800",
  5364 => x"4020",
  5365 => x"F820",
  5366 => x"2020",
  5367 => x"F800",
  5368 => x"5000",
  5369 => x"F820",
  5370 => x"2020",
  5371 => x"F800",
  5372 => x"2050",
  5373 => x"F820",
  5374 => x"2020",
  5375 => x"F800",
  5376 => x"1020",
  5377 => x"7088",
  5378 => x"8888",
  5379 => x"7000",
  5380 => x"4020",
  5381 => x"7088",
  5382 => x"8888",
  5383 => x"7000",
  5384 => x"5000",
  5385 => x"7088",
  5386 => x"8888",
  5387 => x"7000",
  5388 => x"2050",
  5389 => x"7088",
  5390 => x"8888",
  5391 => x"7000",
  5392 => x"1020",
  5393 => x"8888",
  5394 => x"8888",
  5395 => x"7000",
  5396 => x"4020",
  5397 => x"8888",
  5398 => x"8888",
  5399 => x"7000",
  5400 => x"5000",
  5401 => x"8888",
  5402 => x"8888",
  5403 => x"7000",
  5404 => x"2050",
  5405 => x"0088",
  5406 => x"8888",
  5407 => x"7000",
  5408 => x"1020",
  5409 => x"7008",
  5410 => x"7888",
  5411 => x"7800",
  5412 => x"4020",
  5413 => x"7008",
  5414 => x"7888",
  5415 => x"7800",
  5416 => x"5000",
  5417 => x"7008",
  5418 => x"7888",
  5419 => x"7800",
  5420 => x"2050",
  5421 => x"7008",
  5422 => x"7888",
  5423 => x"7800",
  5424 => x"1020",
  5425 => x"7884",
  5426 => x"FC80",
  5427 => x"7C00",
  5428 => x"2010",
  5429 => x"7884",
  5430 => x"FC80",
  5431 => x"7C00",
  5432 => x"5000",
  5433 => x"7884",
  5434 => x"FC80",
  5435 => x"7C00",
  5436 => x"2050",
  5437 => x"7884",
  5438 => x"FC80",
  5439 => x"7C00",
  5440 => x"1020",
  5441 => x"0060",
  5442 => x"2020",
  5443 => x"7000",
  5444 => x"4020",
  5445 => x"0060",
  5446 => x"2020",
  5447 => x"7000",
  5448 => x"0050",
  5449 => x"0060",
  5450 => x"2020",
  5451 => x"7000",
  5452 => x"2050",
  5453 => x"0060",
  5454 => x"2020",
  5455 => x"7000",
  5456 => x"1020",
  5457 => x"0070",
  5458 => x"8888",
  5459 => x"7000",
  5460 => x"4020",
  5461 => x"0070",
  5462 => x"8888",
  5463 => x"7000",
  5464 => x"0050",
  5465 => x"0070",
  5466 => x"8888",
  5467 => x"7000",
  5468 => x"2050",
  5469 => x"0070",
  5470 => x"8888",
  5471 => x"7000",
  5472 => x"1020",
  5473 => x"0088",
  5474 => x"8898",
  5475 => x"6800",
  5476 => x"4020",
  5477 => x"0088",
  5478 => x"8898",
  5479 => x"6800",
  5480 => x"0050",
  5481 => x"0088",
  5482 => x"8898",
  5483 => x"6800",
  5484 => x"2050",
  5485 => x"0088",
  5486 => x"8898",
  5487 => x"6800",
  5488 => x"5000",
  5489 => x"8850",
  5490 => x"2020",
  5491 => x"2000",
  5492 => x"5000",
  5493 => x"8850",
  5494 => x"2040",
  5495 => x"8000",
  5496 => x"2000",
  5497 => x"2040",
  5498 => x"8088",
  5499 => x"7000",
  5500 => x"2020",
  5501 => x"0020",
  5502 => x"2020",
  5503 => x"2000",
  5505 => x"4890",
  5506 => x"4800",
  5509 => x"9048",
  5510 => x"9000",
  5512 => x"8822",
  5513 => x"8822",
  5514 => x"8822",
  5515 => x"8822",
  5516 => x"AA55",
  5517 => x"AA55",
  5518 => x"AA55",
  5519 => x"AA54",
  5520 => x"CCFF",
  5521 => x"33CC",
  5522 => x"FF33",
  5523 => x"CCFF",
  5524 => x"3030",
  5525 => x"3030",
  5526 => x"3030",
  5527 => x"3030",
  5529 => x"00FC",
  5530 => x"FC00",
  5532 => x"3030",
  5533 => x"303C",
  5534 => x"3C00",
  5536 => x"3030",
  5537 => x"30F0",
  5538 => x"F000",
  5541 => x"003C",
  5542 => x"3C30",
  5543 => x"3030",
  5545 => x"00F0",
  5546 => x"F030",
  5547 => x"3030",
  5548 => x"3030",
  5549 => x"30F0",
  5550 => x"F030",
  5551 => x"3030",
  5552 => x"3030",
  5553 => x"30FC",
  5554 => x"FC00",
  5556 => x"3030",
  5557 => x"303C",
  5558 => x"3C30",
  5559 => x"3030",
  5561 => x"00FC",
  5562 => x"FC30",
  5563 => x"3030",
  5564 => x"3030",
  5565 => x"30FC",
  5566 => x"FC30",
  5567 => x"3030",
  5568 => x"3030",
  5569 => x"3030",
  5570 => x"3000",
  5573 => x"00F0",
  5574 => x"F000",
  5577 => x"003C",
  5578 => x"3C00",
  5581 => x"0030",
  5582 => x"3030",
  5583 => x"3030",
  5584 => x"FC84",
  5585 => x"8484",
  5586 => x"8484",
  5587 => x"84FC",
  5588 => x"FCFC",
  5589 => x"CCCC",
  5590 => x"CCCC",
  5591 => x"FCFC",
  5592 => x"FCFC",
  5593 => x"FCFC",
  5594 => x"FCFC",
  5595 => x"FCFC",
  5596 => x"FCFC",
  5597 => x"FCFC",
  5600 => x"E0E0",
  5601 => x"E0E0",
  5602 => x"E0E0",
  5603 => x"E0E0",
  5604 => x"1C1C",
  5605 => x"1C1C",
  5606 => x"1C1C",
  5607 => x"1C1C",
  5610 => x"FCFC",
  5611 => x"FCFC",
  5613 => x"6890",
  5614 => x"9090",
  5615 => x"6800",
  5616 => x"3048",
  5617 => x"4870",
  5618 => x"4868",
  5619 => x"5000",
  5620 => x"00F8",
  5621 => x"8080",
  5622 => x"8080",
  5623 => x"8000",
  5624 => x"0040",
  5625 => x"A810",
  5626 => x"1010",
  5627 => x"1000",
  5628 => x"2020",
  5629 => x"5050",
  5630 => x"8888",
  5631 => x"F800",
  5632 => x"7088",
  5633 => x"6010",
  5634 => x"7088",
  5635 => x"7000",
  5637 => x"7880",
  5638 => x"F880",
  5639 => x"7800",
  5640 => x"2018",
  5641 => x"2040",
  5642 => x"3008",
  5643 => x"7000",
  5644 => x"7088",
  5645 => x"88F8",
  5646 => x"8888",
  5647 => x"7000",
  5649 => x"C040",
  5650 => x"4050",
  5651 => x"2000",
  5652 => x"2020",
  5653 => x"5050",
  5654 => x"8888",
  5655 => x"8800",
  5656 => x"00C0",
  5657 => x"2020",
  5658 => x"5048",
  5659 => x"8800",
  5661 => x"9080",
  5662 => x"90F8",
  5663 => x"8000",
  5664 => x"00F8",
  5665 => x"8888",
  5666 => x"8888",
  5667 => x"8800",
  5669 => x"00F8",
  5670 => x"5050",
  5671 => x"5000",
  5672 => x"FC40",
  5673 => x"2010",
  5674 => x"2040",
  5675 => x"F800",
  5677 => x"7890",
  5678 => x"9090",
  5679 => x"6000",
  5681 => x"78A0",
  5682 => x"2020",
  5683 => x"1800",
  5684 => x"2020",
  5685 => x"70A8",
  5686 => x"7020",
  5687 => x"2000",
  5688 => x"8048",
  5689 => x"5020",
  5690 => x"5090",
  5691 => x"0800",
  5692 => x"0070",
  5693 => x"8888",
  5694 => x"8850",
  5695 => x"D800",
  5696 => x"00F8",
  5697 => x"00F8",
  5698 => x"00F8",
  5700 => x"0020",
  5701 => x"20F8",
  5702 => x"2020",
  5703 => x"F800",
  5704 => x"C030",
  5705 => x"0830",
  5706 => x"C000",
  5707 => x"F800",
  5708 => x"1860",
  5709 => x"8060",
  5710 => x"1800",
  5711 => x"F800",
  5712 => x"0020",
  5713 => x"00F8",
  5714 => x"0020",
  5716 => x"3048",
  5717 => x"3000",
  5720 => x"0018",
  5721 => x"1010",
  5722 => x"9050",
  5723 => x"2000",
  5724 => x"6010",
  5725 => x"2070",
  5728 => x"7088",
  5729 => x"8890",
  5730 => x"8888",
  5731 => x"88B0",
  5732 => x"0020",
  5733 => x"70A0",
  5734 => x"A070",
  5735 => x"2000",
  5736 => x"3C50",
  5737 => x"90FC",
  5738 => x"9090",
  5739 => x"9C00",
  5740 => x"7C90",
  5741 => x"909C",
  5742 => x"9090",
  5743 => x"7C00",
  5744 => x"7088",
  5745 => x"80F0",
  5746 => x"4040",
  5747 => x"F800",
  5748 => x"8888",
  5749 => x"50F8",
  5750 => x"20F8",
  5751 => x"2000",
  5752 => x"1028",
  5753 => x"2020",
  5754 => x"20A0",
  5755 => x"4000",
  5756 => x"F880",
  5757 => x"80F0",
  5758 => x"8888",
  5759 => x"F000",
  5760 => x"F050",
  5761 => x"5090",
  5762 => x"90F8",
  5763 => x"8800",
  5764 => x"A8A8",
  5765 => x"70A8",
  5766 => x"A8A8",
  5767 => x"A800",
  5768 => x"7088",
  5769 => x"0830",
  5770 => x"0888",
  5771 => x"7000",
  5772 => x"8888",
  5773 => x"C8A8",
  5774 => x"9888",
  5775 => x"8800",
  5776 => x"5020",
  5777 => x"88C8",
  5778 => x"A898",
  5779 => x"8800",
  5780 => x"7848",
  5781 => x"4848",
  5782 => x"4848",
  5783 => x"C800",
  5784 => x"8888",
  5785 => x"8888",
  5786 => x"88F8",
  5787 => x"0800",
  5788 => x"8888",
  5789 => x"8878",
  5790 => x"0808",
  5791 => x"0800",
  5792 => x"A8A8",
  5793 => x"A8A8",
  5794 => x"A8A8",
  5795 => x"F800",
  5796 => x"A8A8",
  5797 => x"A8A8",
  5798 => x"A8F8",
  5799 => x"0800",
  5800 => x"C040",
  5801 => x"4070",
  5802 => x"4848",
  5803 => x"7000",
  5804 => x"8888",
  5805 => x"88E8",
  5806 => x"9898",
  5807 => x"E800",
  5808 => x"8080",
  5809 => x"80F0",
  5810 => x"8888",
  5811 => x"F000",
  5812 => x"7088",
  5813 => x"0878",
  5814 => x"0888",
  5815 => x"7000",
  5816 => x"90A8",
  5817 => x"A8E8",
  5818 => x"A8A8",
  5819 => x"9000",
  5820 => x"7888",
  5821 => x"8878",
  5822 => x"4888",
  5823 => x"8800",
  5824 => x"4865",
  5825 => x"6C6C",
  5826 => x"6F20",
  5827 => x"576F",
  5828 => x"726C",
  5829 => x"643F",
  5830 => x"0041",
  5831 => x"6E6F",
  5832 => x"7468",
  5833 => x"6572",
  5834 => x"2074",
  5835 => x"6573",
  5836 => x"7400",
  others => x"0000"
 );
begin
   process(CLK)
	begin 
		if (CLK'event AND CLK='1') then
			DOUT2 <= memoire(to_integer(unsigned(AD2)));
		end if;
	end process;

	process(CLK)
	begin 
		if (CLK'event AND CLK='1') then
			if ((CE1='1') AND (OE1='1')) then 
				DOUT1<=memoire(to_integer(unsigned(AD1)));
			else 
				DOUT1<=(others =>'0');
			end if;		
		end if;
	end process;
	
	process (CLK)
	begin
	  IF (CLK'event AND CLK='1') then
			if ((CE1='1') AND (WE1='1')) then 
				memoire(to_integer(unsigned(AD1)))<=DIN1;
			end if;
		  end if;
	end process;
	
end Behavioral;
