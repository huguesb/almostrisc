----------------------------------------------------------------------------------
--
-- File retrieved, on 07/02/2010, from :
-- http://sebastien-viardot.imag.fr/Enseignements/Archi1A2s/sources/ROMPROG.vhd
--
-- Slightly altered to get rid of vendor-specific packages and adjust formatting
-- Now auto-filled by asrom script
--
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROMPROG is
  Port ( AD : in  STD_LOGIC_VECTOR (12 downto 0);
         D : out  STD_LOGIC_VECTOR (15 downto 0);
         CLK : in STD_LOGIC);
end ROMPROG;

architecture Behavioral of ROMPROG is
  constant low_address: natural := 0;
  constant high_address: natural := 8192;
  subtype octet is std_logic_vector( 15 downto 0 );
  type zone_memoire is
    array (natural range low_address to high_address-1) of octet;
  constant m: zone_memoire:= (
    0=>x"FFF7",	-- 1111111111110111  liw	r7, IRQ_mask
    1=>x"2000",	-- 0010000000000000  
    2=>x"F8C0",	-- 1111100011000000  bai	-, os_init
    3=>x"0100",	-- 0000000100000000  
   16=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_ack
   17=>x"2002",	-- 0010000000000010  
   18=>x"D001",	-- 1101000000000001  lw	r1, r0
   19=>x"F54A",	-- 1111010101001010  bspl	r2, r1, 5
   20=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_error
   21=>x"0050",	-- 0000000001010000  
   22=>x"F4CA",	-- 1111010011001010  bspl	r2, r1, 3
   23=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_kbd
   24=>x"0060",	-- 0000000001100000  
   25=>x"F40A",	-- 1111010000001010  bspl	r2, r1, 0
   26=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_tmr
   27=>x"0040",	-- 0000000001000000  
   28=>x"D201",	-- 1101001000000001  sw	r1, r0
   29=>x"FFFE",	-- 1111111111111110  reti
   64=>x"263F",	-- 0010011000111111  not r7, r7
   65=>x"D7C0",	-- 1101011111000000  out	r7
   66=>x"E383",	-- 1110001110000011  ba	-, r6
   80=>x"25FF",	-- 0010010111111111  xor	r7, r7, r7
   81=>x"D7C0",	-- 1101011111000000  out	r7
   82=>x"E383",	-- 1110001110000011  ba	-, r6
   96=>x"FFF2",	-- 1111111111110010  liw	r2, PS2_rx
   97=>x"2004",	-- 0010000000000100  
   98=>x"D012",	-- 1101000000010010  lw	r2, r2
   99=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map + 8
  100=>x"16C8",	-- 0001011011001000  
  101=>x"D01B",	-- 1101000000011011  lw	r3, r3
  102=>x"1EBF",	-- 0001111010111111  mixll	r7, r7, r2
  103=>x"C784",	-- 1100011110000100  li	r4, 0xF0
  104=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  105=>x"8B20",	-- 1000101100100000  brieq	r4, int_kbd.release
  106=>x"C704",	-- 1100011100000100  li	r4, 0xE0
  107=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  108=>x"88E0",	-- 1000100011100000  brieq	r4, int_kbd.extended
  109=>x"FFF5",	-- 1111111111110101  liw	r5, paper_keys - 1
  110=>x"16CF",	-- 0001011011001111  
  111=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  112=>x"80E0",	-- 1000000011100000  brieq	r4, $+3
  113=>x"FFF5",	-- 1111111111110101  liw	r5, paper_keys + 11 - 1
  114=>x"16DA",	-- 0001011011011010  
  115=>x"042D",	-- 0000010000101101  inc	r5, r5
  116=>x"D02C",	-- 1101000000101100  lw	r4, r5
  117=>x"8560",	-- 1000010101100000  brieq	r4, scan_code_mismatch
  118=>x"6E24",	-- 0110111000100100  shr	r4, r4, 7
  119=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  120=>x"BEE4",	-- 1011111011100100  brine	r4, scan_code_loop
  121=>x"D02A",	-- 1101000000101010  lw	r2, r5
  122=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  123=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  124=>x"741B",	-- 0111010000011011  shr	r3, r3, 10
  125=>x"C00D",	-- 1100000000001101  li	r5, 1
  126=>x"0612",	-- 0000011000010010  dec	r2, r2
  127=>x"3AAA",	-- 0011101010101010  rrl	r2, r5, r2
  128=>x"FFF5",	-- 1111111111110101  liw	r5, key_press_map
  129=>x"16C0",	-- 0001011011000000  
  130=>x"08ED",	-- 0000100011101101  add	r5, r5, r3
  131=>x"D02B",	-- 1101000000101011  lw	r3, r5
  132=>x"80E4",	-- 1000000011100100  brine	r4, scan_code_release
  133=>x"229B",	-- 0010001010011011  or	r3, r3, r2
  134=>x"80C3",	-- 1000000011000011  bri	-, scan_code_notify
  135=>x"2612",	-- 0010011000010010  not	r2, r2
  136=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  137=>x"D22B",	-- 1101001000101011  sw	r3, r5
  138=>x"C003",	-- 1100000000000011  li	r3, 0
  139=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  140=>x"16C8",	-- 0001011011001000  
  141=>x"D223",	-- 1101001000100011  sw	r3, r4
  142=>x"E383",	-- 1110001110000011  ba	-, r6
  143=>x"C014",	-- 1100000000010100  li	r4, 2
  144=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  145=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  146=>x"16C8",	-- 0001011011001000  
  147=>x"D223",	-- 1101001000100011  sw	r3, r4
  148=>x"E383",	-- 1110001110000011  ba	-, r6
  149=>x"C00C",	-- 1100000000001100  li	r4, 1
  150=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  151=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  152=>x"16C8",	-- 0001011011001000  
  153=>x"D223",	-- 1101001000100011  sw	r3, r4
  154=>x"E383",	-- 1110001110000011  ba	-, r6
  256=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_mask
  257=>x"2000",	-- 0010000000000000  
  258=>x"C0C9",	-- 1100000011001001  li	r1, 0x19
  259=>x"D201",	-- 1101001000000001  sw	r1, r0
  260=>x"0400",	-- 0000010000000000  inc	r0, r0
  261=>x"CFF9",	-- 1100111111111001  li	r1, -1
  262=>x"D201",	-- 1101001000000001  sw	r1, r0
  263=>x"C03A",	-- 1100000000111010  li	r2, 7
  264=>x"0880",	-- 0000100010000000  add	r0, r0, r2
  265=>x"C0EA",	-- 1100000011101010  li	r2, 0x1D
  266=>x"D202",	-- 1101001000000010  sw	r2, r0
  267=>x"0400",	-- 0000010000000000  inc	r0, r0
  268=>x"C07A",	-- 1100000001111010  li	r2, 15
  269=>x"D202",	-- 1101001000000010  sw	r2, r0
  270=>x"0400",	-- 0000010000000000  inc	r0, r0
  271=>x"C0DA",	-- 1100000011011010  li	r2, 0x1B
  272=>x"D202",	-- 1101001000000010  sw	r2, r0
  273=>x"0400",	-- 0000010000000000  inc	r0, r0
  274=>x"FFF2",	-- 1111111111110010  liw	r2, 817
  275=>x"0331",	-- 0000001100110001  
  276=>x"D202",	-- 1101001000000010  sw	r2, r0
  277=>x"FFF0",	-- 1111111111110000  liw	r0, key_press_map
  278=>x"16C0",	-- 0001011011000000  
  279=>x"C001",	-- 1100000000000001  li	r1, 0
  280=>x"C042",	-- 1100000001000010  li	r2, 8
  281=>x"D201",	-- 1101001000000001  sw	r1, r0
  282=>x"0400",	-- 0000010000000000  inc	r0, r0
  283=>x"0612",	-- 0000011000010010  dec	r2, r2
  284=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  285=>x"C0F3",	-- 1100000011110011  li	r3, 30
  286=>x"CFFA",	-- 1100111111111010  li	r2, -1
  287=>x"D21A",	-- 1101001000011010  sw	r2, r3
  288=>x"8083",	-- 1000000010000011  bri	-, PaperGameStart
  289=>x"8003",	-- 1000000000000011  bri	-, PaperMenuLoop
  290=>x"FFF0",	-- 1111111111110000  liw	r0, paper_dir
  291=>x"179C",	-- 0001011110011100  
  292=>x"C001",	-- 1100000000000001  li	r1, 0
  293=>x"D201",	-- 1101001000000001  sw	r1, r0
  294=>x"0400",	-- 0000010000000000  inc	r0, r0
  295=>x"FFF1",	-- 1111111111110001  liw	r1, 152 * 8
  296=>x"04C0",	-- 0000010011000000  
  297=>x"D201",	-- 1101001000000001  sw	r1, r0
  298=>x"0400",	-- 0000010000000000  inc	r0, r0
  299=>x"C001",	-- 1100000000000001  li	r1, 0
  300=>x"D201",	-- 1101001000000001  sw	r1, r0
  301=>x"0400",	-- 0000010000000000  inc	r0, r0
  302=>x"FFF1",	-- 1111111111110001  liw	r1, 128 * 8
  303=>x"0400",	-- 0000010000000000  
  304=>x"D201",	-- 1101001000000001  sw	r1, r0
  305=>x"0400",	-- 0000010000000000  inc	r0, r0
  306=>x"C001",	-- 1100000000000001  li	r1, 0
  307=>x"D201",	-- 1101001000000001  sw	r1, r0
  308=>x"0400",	-- 0000010000000000  inc	r0, r0
  309=>x"C029",	-- 1100000000101001  li	r1, 5
  310=>x"D201",	-- 1101001000000001  sw	r1, r0
  311=>x"0400",	-- 0000010000000000  inc	r0, r0
  312=>x"C011",	-- 1100000000010001  li	r1, 2
  313=>x"D201",	-- 1101001000000001  sw	r1, r0
  314=>x"0400",	-- 0000010000000000  inc	r0, r0
  315=>x"FFF0",	-- 1111111111110000  liw	r0, TMR_cur1
  316=>x"200D",	-- 0010000000001101  
  317=>x"D000",	-- 1101000000000000  lw	r0, r0
  318=>x"FAC6",	-- 1111101011000110  bail	-, r6, rand16_init
  319=>x"0226",	-- 0000001000100110  
  320=>x"C000",	-- 1100000000000000  li	r0, 0
  321=>x"CFF9",	-- 1100111111111001  li	r1, -1
  322=>x"C0A2",	-- 1100000010100010  li	r2, 20
  323=>x"D201",	-- 1101001000000001  sw	r1, r0
  324=>x"0400",	-- 0000010000000000  inc	r0, r0
  325=>x"0612",	-- 0000011000010010  dec	r2, r2
  326=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  327=>x"C001",	-- 1100000000000001  li	r1, 0
  328=>x"FFF2",	-- 1111111111110010  liw	r2, 18*20
  329=>x"0168",	-- 0000000101101000  
  330=>x"D201",	-- 1101001000000001  sw	r1, r0
  331=>x"0400",	-- 0000010000000000  inc	r0, r0
  332=>x"0612",	-- 0000011000010010  dec	r2, r2
  333=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  334=>x"CFF9",	-- 1100111111111001  li	r1, -1
  335=>x"C0A2",	-- 1100000010100010  li	r2, 20
  336=>x"D201",	-- 1101001000000001  sw	r1, r0
  337=>x"0400",	-- 0000010000000000  inc	r0, r0
  338=>x"0612",	-- 0000011000010010  dec	r2, r2
  339=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  340=>x"C020",	-- 1100000000100000  li	r0, 4
  341=>x"C029",	-- 1100000000101001  li	r1, 5
  342=>x"FFF2",	-- 1111111111110010  liw	r2, paper_title
  343=>x"17A4",	-- 0001011110100100  
  344=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  345=>x"026C",	-- 0000001001101100  
  346=>x"C778",	-- 1100011101111000  li	r0, 239
  347=>x"C009",	-- 1100000000001001  li	r1, 1
  348=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud
  349=>x"1780",	-- 0001011110000000  
  350=>x"C043",	-- 1100000001000011  li	r3, 8
  351=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  352=>x"036E",	-- 0000001101101110  
  353=>x"C0F8",	-- 1100000011111000  li	r0, 31
  354=>x"C009",	-- 1100000000001001  li	r1, 1
  355=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed + 1
  356=>x"17A1",	-- 0001011110100001  
  357=>x"D012",	-- 1101000000010010  lw	r2, r2
  358=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum
  359=>x"029B",	-- 0000001010011011  
  360=>x"C120",	-- 1100000100100000  li	r0, 36
  361=>x"C009",	-- 1100000000001001  li	r1, 1
  362=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  363=>x"17AA",	-- 0001011110101010  
  364=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  365=>x"026C",	-- 0000001001101100  
  366=>x"C778",	-- 1100011101111000  li	r0, 239
  367=>x"C051",	-- 1100000001010001  li	r1, 10
  368=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud + 4
  369=>x"1784",	-- 0001011110000100  
  370=>x"C043",	-- 1100000001000011  li	r3, 8
  371=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  372=>x"036E",	-- 0000001101101110  
  373=>x"C0F8",	-- 1100000011111000  li	r0, 31
  374=>x"C051",	-- 1100000001010001  li	r1, 10
  375=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed + 2
  376=>x"17A2",	-- 0001011110100010  
  377=>x"D012",	-- 1101000000010010  lw	r2, r2
  378=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum
  379=>x"029B",	-- 0000001010011011  
  380=>x"C120",	-- 1100000100100000  li	r0, 36
  381=>x"C051",	-- 1100000001010001  li	r1, 10
  382=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  383=>x"17AA",	-- 0001011110101010  
  384=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  385=>x"026C",	-- 0000001001101100  
  386=>x"FFF0",	-- 1111111111110000  liw	r0, 20*20
  387=>x"0190",	-- 0000000110010000  
  388=>x"C001",	-- 1100000000000001  li	r1, 0
  389=>x"FFF2",	-- 1111111111110010  liw	r2, 220*20
  390=>x"1130",	-- 0001000100110000  
  391=>x"D201",	-- 1101001000000001  sw	r1, r0
  392=>x"0400",	-- 0000010000000000  inc	r0, r0
  393=>x"0612",	-- 0000011000010010  dec	r2, r2
  394=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  395=>x"FFF5",	-- 1111111111110101  liw	r5, paper_tilemap
  396=>x"17B0",	-- 0001011110110000  
  397=>x"D02C",	-- 1101000000101100  lw	r4, r5
  398=>x"042D",	-- 0000010000101101  inc	r5, r5
  399=>x"88E0",	-- 1000100011100000  brieq	r4, PaperGameTileSkip
  400=>x"063F",	-- 0000011000111111  dec	r7, r7
  401=>x"D23D",	-- 1101001000111101  sw	r5, r7
  402=>x"FFF3",	-- 1111111111110011  liw	r3, paper_tilemap
  403=>x"17B0",	-- 0001011110110000  
  404=>x"0AEB",	-- 0000101011101011  sub	r3, r5, r3
  405=>x"6E20",	-- 0110111000100000  shr	r0, r4, 7
  406=>x"6219",	-- 0110001000011001  shr	r1, r3, 1
  407=>x"4409",	-- 0100010000001001  shl	r1, r1, 2
  408=>x"C0DA",	-- 1100000011011010  li	r2, 27
  409=>x"0889",	-- 0000100010001001  add	r1, r1, r2
  410=>x"FFF2",	-- 1111111111110010  liw	r2, paper_pos + 1
  411=>x"179E",	-- 0001011110011110  
  412=>x"D012",	-- 1101000000010010  lw	r2, r2
  413=>x"6412",	-- 0110010000010010  shr	r2, r2, 2
  414=>x"C03B",	-- 1100000000111011  li	r3, 7
  415=>x"20D2",	-- 0010000011010010  and	r2, r2, r3
  416=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  417=>x"4E24",	-- 0100111000100100  shl	r4, r4, 7
  418=>x"6E24",	-- 0110111000100100  shr	r4, r4, 7
  419=>x"C00B",	-- 1100000000001011  li	r3, 1
  420=>x"FB06",	-- 1111101100000110  bailne	r0, r6, put_tile
  421=>x"023C",	-- 0000001000111100  
  422=>x"C013",	-- 1100000000010011  li	r3, 2
  423=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_tile
  424=>x"023C",	-- 0000001000111100  
  425=>x"0624",	-- 0000011000100100  dec	r4, r4
  426=>x"BF64",	-- 1011111101100100  brine	r4, PaperGameSegmentLoop
  427=>x"C003",	-- 1100000000000011  li	r3, 0
  428=>x"C144",	-- 1100000101000100  li	r4, 40
  429=>x"0B04",	-- 0000101100000100  sub	r4, r0, r4
  430=>x"FB66",	-- 1111101101100110  baillt	r4, r6, put_tile
  431=>x"023C",	-- 0000001000111100  
  432=>x"D03D",	-- 1101000000111101  lw	r5, r7
  433=>x"043F",	-- 0000010000111111  inc	r7, r7
  434=>x"FFF4",	-- 1111111111110100  liw r4, paper_tilemap + 125
  435=>x"182D",	-- 0001100000101101  
  436=>x"0B2C",	-- 0000101100101100  sub	r4, r5, r4
  437=>x"B625",	-- 1011011000100101  brilt	r4, PaperGameTileLoop
  438=>x"FFF3",	-- 1111111111110011  liw	r3, paper_speed
  439=>x"17A0",	-- 0001011110100000  
  440=>x"D01B",	-- 1101000000011011  lw	r3, r3
  441=>x"CFC4",	-- 1100111111000100  li	r4, 0x1F8
  442=>x"211C",	-- 0010000100011100  and	r4, r3, r4
  443=>x"0924",	-- 0000100100100100  add	r4, r4, r4
  444=>x"0924",	-- 0000100100100100  add	r4, r4, r4
  445=>x"FFF3",	-- 1111111111110011  liw	r3, paper_pos
  446=>x"179D",	-- 0001011110011101  
  447=>x"D018",	-- 1101000000011000  lw	r0, r3
  448=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  449=>x"FFF2",	-- 1111111111110010  liw	r2, paper_sprites
  450=>x"1720",	-- 0001011100100000  
  451=>x"0912",	-- 0000100100010010  add	r2, r2, r4
  452=>x"C161",	-- 1100000101100001  li	r1, 44
  453=>x"C083",	-- 1100000010000011  li	r3, 16
  454=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_16_masked
  455=>x"0308",	-- 0000001100001000  
  456=>x"942C",	-- 1001010000101100  brine	r5, PaperGameFail
  458=>x"C028",	-- 1100000000101000  li	r0, 5
  459=>x"C001",	-- 1100000000000001  li	r1, 0
  460=>x"8043",	-- 1000000001000011  bri	-, $+1
  461=>x"8043",	-- 1000000001000011  bri	-, $+1
  462=>x"0609",	-- 0000011000001001  dec	r1, r1
  463=>x"BF4C",	-- 1011111101001100  brine	r1, $-3
  464=>x"0600",	-- 0000011000000000  dec	r0, r0
  465=>x"BE84",	-- 1011111010000100  brine	r0, $-6
  466=>x"FFF2",	-- 1111111111110010  liw	r2, paper_pos
  467=>x"179D",	-- 0001011110011101  
  468=>x"FFF3",	-- 1111111111110011  liw	r3, paper_speed
  469=>x"17A0",	-- 0001011110100000  
  470=>x"D010",	-- 1101000000010000  lw	r0, r2
  471=>x"D019",	-- 1101000000011001  lw	r1, r3
  472=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  473=>x"8FC5",	-- 1000111111000101  brilt	r0, PaperGameFail
  474=>x"FFF4",	-- 1111111111110100  liw	r4, 304*8
  475=>x"0980",	-- 0000100110000000  
  476=>x"0B04",	-- 0000101100000100  sub	r4, r0, r4
  477=>x"8EE1",	-- 1000111011100001  brige	r4, PaperGameFail
  478=>x"D210",	-- 1101001000010000  sw	r0, r2
  479=>x"0412",	-- 0000010000010010  inc	r2, r2
  480=>x"041B",	-- 0000010000011011  inc	r3, r3
  481=>x"D010",	-- 1101000000010000  lw	r0, r2
  482=>x"D019",	-- 1101000000011001  lw	r1, r3
  483=>x"C1FC",	-- 1100000111111100  li	r4, 0x3F
  484=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  485=>x"2101",	-- 0010000100000001  and	r1, r0, r4
  486=>x"2624",	-- 0010011000100100  not	r4, r4
  487=>x"2100",	-- 0010000100000000  and	r0, r0, r4
  488=>x"D211",	-- 1101001000010001  sw	r1, r2
  489=>x"8480",	-- 1000010010000000  brieq	r0, PaperGameSkipScroll
  490=>x"FFF0",	-- 1111111111110000  liw	r0, paper_tilemap
  491=>x"17B0",	-- 0001011110110000  
  492=>x"C021",	-- 1100000000100001  li	r1, 4
  493=>x"0841",	-- 0000100001000001  add	r1, r0, r1
  494=>x"C302",	-- 1100001100000010  li	r2, 24*4
  495=>x"D00B",	-- 1101000000001011  lw	r3, r1
  496=>x"D203",	-- 1101001000000011  sw	r3, r0
  497=>x"0400",	-- 0000010000000000  inc	r0, r0
  498=>x"0409",	-- 0000010000001001  inc	r1, r1
  499=>x"0612",	-- 0000011000010010  dec	r2, r2
  500=>x"BED4",	-- 1011111011010100  brine	r2, PaperGameScrollLoop
  501=>x"C03A",	-- 1100000000111010  li	r2, 7
  502=>x"640B",	-- 0110010000001011  shr	r3, r1, 2
  503=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  504=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  505=>x"1EC9",	-- 0001111011001001  mixll	r1, r1, r3
  506=>x"D201",	-- 1101001000000001  sw	r1, r0
  507=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  508=>x"16C0",	-- 0001011011000000  
  509=>x"D01B",	-- 1101000000011011  lw	r3, r3
  510=>x"F818",	-- 1111100000011000  baieq	r3, PaperGameRedrawContent
  511=>x"0182",	-- 0000000110000010  
  512=>x"F7DC",	-- 1111011111011100  bspl	r4, r3, 15
  513=>x"8924",	-- 1000100100100100  brine	r4, PaperGameQuit
  514=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  515=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveUp
  516=>x"F49C",	-- 1111010010011100  bspl	r4, r3, 2
  517=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveDOWN
  518=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  519=>x"81E0",	-- 1000000111100000  brieq	r4, PaperNoMoveLEFT
  520=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  521=>x"17A0",	-- 0001011110100000  
  522=>x"D010",	-- 1101000000010000  lw	r0, r2
  523=>x"0600",	-- 0000011000000000  dec	r0, r0
  524=>x"0600",	-- 0000011000000000  dec	r0, r0
  525=>x"D210",	-- 1101001000010000  sw	r0, r2
  526=>x"F4DC",	-- 1111010011011100  bspl	r4, r3, 3
  527=>x"81E0",	-- 1000000111100000  brieq	r4, PaperNoMoveRIGHT
  528=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  529=>x"17A0",	-- 0001011110100000  
  530=>x"D010",	-- 1101000000010000  lw	r0, r2
  531=>x"0400",	-- 0000010000000000  inc	r0, r0
  532=>x"0400",	-- 0000010000000000  inc	r0, r0
  533=>x"D210",	-- 1101001000010000  sw	r0, r2
  534=>x"F8C0",	-- 1111100011000000  bai	-, PaperGameRedrawContent
  535=>x"0182",	-- 0000000110000010  
  536=>x"C000",	-- 1100000000000000  li	r0, 0
  537=>x"FFF2",	-- 1111111111110010  liw	r2, 240*20
  538=>x"12C0",	-- 0001001011000000  
  539=>x"D001",	-- 1101000000000001  lw	r1, r0
  540=>x"2609",	-- 0010011000001001  not	r1, r1
  541=>x"D201",	-- 1101001000000001  sw	r1, r0
  542=>x"0400",	-- 0000010000000000  inc	r0, r0
  543=>x"0612",	-- 0000011000010010  dec	r2, r2
  544=>x"BED4",	-- 1011111011010100  brine	r2, $-5
  545=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  546=>x"16C0",	-- 0001011011000000  
  547=>x"D01A",	-- 1101000000011010  lw	r2, r3
  548=>x"BFD0",	-- 1011111111010000  brieq	r2, $-1
  549=>x"FFFF",	-- 1111111111111111  reset
  550=>x"FFF2",	-- 1111111111110010  liw	r2, rand_seed
  551=>x"16C8",	-- 0001011011001000  
  552=>x"D210",	-- 1101001000010000  sw	r0, r2
  553=>x"E383",	-- 1110001110000011  ba	-, r6
  554=>x"FFF2",	-- 1111111111110010  liw	r2, rand_seed
  555=>x"16C8",	-- 0001011011001000  
  556=>x"D013",	-- 1101000000010011  lw	r3, r2
  557=>x"C7EC",	-- 1100011111101100  li	r4, 253
  558=>x"1F19",	-- 0001111100011001  mixll	r1, r3, r4
  559=>x"18E4",	-- 0001100011100100  mixhh	r4, r4, r3
  560=>x"C002",	-- 1100000000000010  li	r2, 0
  561=>x"0AC9",	-- 0000101011001001  sub	r1, r1, r3
  562=>x"0EA4",	-- 0000111010100100  sbc	r4, r4, r2
  563=>x"0EC9",	-- 0000111011001001  sbc	r1, r1, r3
  564=>x"0EA4",	-- 0000111010100100  sbc	r4, r4, r2
  565=>x"1B13",	-- 0001101100010011  mixhl	r3, r2, r4
  566=>x"0EC9",	-- 0000111011001001  sbc	r1, r1, r3
  567=>x"0C89",	-- 0000110010001001  adc	r1, r1, r2
  568=>x"FFF2",	-- 1111111111110010  liw	r2, rand_seed
  569=>x"16C8",	-- 0001011011001000  
  570=>x"D211",	-- 1101001000010001  sw	r1, r2
  571=>x"E383",	-- 1110001110000011  ba	-, r6
  572=>x"063F",	-- 0000011000111111  dec	r7, r7
  573=>x"D238",	-- 1101001000111000  sw	r0, r7
  574=>x"063F",	-- 0000011000111111  dec	r7, r7
  575=>x"D239",	-- 1101001000111001  sw	r1, r7
  576=>x"063F",	-- 0000011000111111  dec	r7, r7
  577=>x"D23A",	-- 1101001000111010  sw	r2, r7
  578=>x"063F",	-- 0000011000111111  dec	r7, r7
  579=>x"D23B",	-- 1101001000111011  sw	r3, r7
  580=>x"063F",	-- 0000011000111111  dec	r7, r7
  581=>x"D23C",	-- 1101001000111100  sw	r4, r7
  582=>x"063F",	-- 0000011000111111  dec	r7, r7
  583=>x"D23D",	-- 1101001000111101  sw	r5, r7
  584=>x"063F",	-- 0000011000111111  dec	r7, r7
  585=>x"D23E",	-- 1101001000111110  sw	r6, r7
  586=>x"FFF2",	-- 1111111111110010  liw	r2, paper_tiles
  587=>x"1790",	-- 0001011110010000  
  588=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  589=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  590=>x"C043",	-- 1100000001000011  li	r3, 8
  591=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  592=>x"0348",	-- 0000001101001000  
  593=>x"D03E",	-- 1101000000111110  lw	r6, r7
  594=>x"043F",	-- 0000010000111111  inc	r7, r7
  595=>x"D03D",	-- 1101000000111101  lw	r5, r7
  596=>x"043F",	-- 0000010000111111  inc	r7, r7
  597=>x"D03C",	-- 1101000000111100  lw	r4, r7
  598=>x"043F",	-- 0000010000111111  inc	r7, r7
  599=>x"D03B",	-- 1101000000111011  lw	r3, r7
  600=>x"043F",	-- 0000010000111111  inc	r7, r7
  601=>x"D03A",	-- 1101000000111010  lw	r2, r7
  602=>x"043F",	-- 0000010000111111  inc	r7, r7
  603=>x"D039",	-- 1101000000111001  lw	r1, r7
  604=>x"043F",	-- 0000010000111111  inc	r7, r7
  605=>x"D038",	-- 1101000000111000  lw	r0, r7
  606=>x"043F",	-- 0000010000111111  inc	r7, r7
  607=>x"0400",	-- 0000010000000000  inc	r0, r0
  608=>x"E383",	-- 1110001110000011  ba	-, r6
  609=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  610=>x"C084",	-- 1100000010000100  li	r4, 16
  611=>x"0800",	-- 0000100000000000  add	r0, r0, r0
  612=>x"0C49",	-- 0000110001001001  adc	r1, r1, r1
  613=>x"0A8B",	-- 0000101010001011  sub	r3, r1, r2
  614=>x"80DD",	-- 1000000011011101  brilt	r3, div_16_16.skip
  615=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  616=>x"0400",	-- 0000010000000000  inc	r0, r0
  617=>x"0624",	-- 0000011000100100  dec	r4, r4
  618=>x"BE64",	-- 1011111001100100  brine	r4, div_16_16.loop
  619=>x"E383",	-- 1110001110000011  ba	-, r6
  620=>x"063F",	-- 0000011000111111  dec	r7, r7
  621=>x"D23E",	-- 1101001000111110  sw	r6, r7
  622=>x"D013",	-- 1101000000010011  lw	r3, r2
  623=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  624=>x"84D8",	-- 1000010011011000  brieq	r3, puts.end
  625=>x"063F",	-- 0000011000111111  dec	r7, r7
  626=>x"D23A",	-- 1101001000111010  sw	r2, r7
  627=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  628=>x"0286",	-- 0000001010000110  
  629=>x"D03A",	-- 1101000000111010  lw	r2, r7
  630=>x"043F",	-- 0000010000111111  inc	r7, r7
  631=>x"D013",	-- 1101000000010011  lw	r3, r2
  632=>x"4E1B",	-- 0100111000011011  shl	r3, r3, 7
  633=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  634=>x"8258",	-- 1000001001011000  brieq	r3, puts.end
  635=>x"063F",	-- 0000011000111111  dec	r7, r7
  636=>x"D23A",	-- 1101001000111010  sw	r2, r7
  637=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  638=>x"0286",	-- 0000001010000110  
  639=>x"D03A",	-- 1101000000111010  lw	r2, r7
  640=>x"043F",	-- 0000010000111111  inc	r7, r7
  641=>x"0412",	-- 0000010000010010  inc	r2, r2
  642=>x"BB03",	-- 1011101100000011  bri	-, puts.loop
  643=>x"D03E",	-- 1101000000111110  lw	r6, r7
  644=>x"043F",	-- 0000010000111111  inc	r7, r7
  645=>x"E383",	-- 1110001110000011  ba	-, r6
  646=>x"063F",	-- 0000011000111111  dec	r7, r7
  647=>x"D23E",	-- 1101001000111110  sw	r6, r7
  648=>x"063F",	-- 0000011000111111  dec	r7, r7
  649=>x"D238",	-- 1101001000111000  sw	r0, r7
  650=>x"063F",	-- 0000011000111111  dec	r7, r7
  651=>x"D239",	-- 1101001000111001  sw	r1, r7
  652=>x"FFF2",	-- 1111111111110010  liw	r2, font_map
  653=>x"12C0",	-- 0001001011000000  
  654=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  655=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  656=>x"C043",	-- 1100000001000011  li	r3, 8
  657=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  658=>x"0348",	-- 0000001101001000  
  659=>x"D039",	-- 1101000000111001  lw	r1, r7
  660=>x"043F",	-- 0000010000111111  inc	r7, r7
  661=>x"D038",	-- 1101000000111000  lw	r0, r7
  662=>x"043F",	-- 0000010000111111  inc	r7, r7
  663=>x"0400",	-- 0000010000000000  inc	r0, r0
  664=>x"D03E",	-- 1101000000111110  lw	r6, r7
  665=>x"043F",	-- 0000010000111111  inc	r7, r7
  666=>x"E383",	-- 1110001110000011  ba	-, r6
  667=>x"063F",	-- 0000011000111111  dec	r7, r7
  668=>x"D23E",	-- 1101001000111110  sw	r6, r7
  669=>x"FFF4",	-- 1111111111110100  liw	r4, 10000
  670=>x"2710",	-- 0010011100010000  
  671=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  672=>x"02AE",	-- 0000001010101110  
  673=>x"FFF4",	-- 1111111111110100  liw	r4, 1000
  674=>x"03E8",	-- 0000001111101000  
  675=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  676=>x"02AE",	-- 0000001010101110  
  677=>x"C324",	-- 1100001100100100  li	r4, 100
  678=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  679=>x"02AE",	-- 0000001010101110  
  680=>x"C054",	-- 1100000001010100  li	r4, 10
  681=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  682=>x"02AE",	-- 0000001010101110  
  683=>x"D03E",	-- 1101000000111110  lw	r6, r7
  684=>x"043F",	-- 0000010000111111  inc	r7, r7
  685=>x"C00C",	-- 1100000000001100  li	r4, 1
  686=>x"C17B",	-- 1100000101111011  li	r3, 0x2F
  687=>x"041B",	-- 0000010000011011  inc	r3, r3
  688=>x"0B12",	-- 0000101100010010  sub	r2, r2, r4
  689=>x"BF91",	-- 1011111110010001  brige	r2, printnum.loop
  690=>x"0912",	-- 0000100100010010  add	r2, r2, r4
  691=>x"063F",	-- 0000011000111111  dec	r7, r7
  692=>x"D23E",	-- 1101001000111110  sw	r6, r7
  693=>x"063F",	-- 0000011000111111  dec	r7, r7
  694=>x"D23A",	-- 1101001000111010  sw	r2, r7
  695=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  696=>x"0286",	-- 0000001010000110  
  697=>x"D03A",	-- 1101000000111010  lw	r2, r7
  698=>x"043F",	-- 0000010000111111  inc	r7, r7
  699=>x"D03E",	-- 1101000000111110  lw	r6, r7
  700=>x"043F",	-- 0000010000111111  inc	r7, r7
  701=>x"E383",	-- 1110001110000011  ba	-, r6
  702=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  703=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  704=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  705=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  706=>x"C0A0",	-- 1100000010100000  li	r0, 20
  707=>x"0412",	-- 0000010000010010  inc	r2, r2
  708=>x"D011",	-- 1101000000010001  lw	r1, r2
  709=>x"E421",	-- 1110010000100001  exw	r1, r4
  710=>x"0412",	-- 0000010000010010  inc	r2, r2
  711=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  712=>x"061B",	-- 0000011000011011  dec	r3, r3
  713=>x"BE9C",	-- 1011111010011100  brine	r3, put_sprite_16_aligned.loop
  714=>x"C005",	-- 1100000000000101  li	r5, 0
  715=>x"E383",	-- 1110001110000011  ba	-, r6
  716=>x"C07D",	-- 1100000001111101  li	r5, 15
  717=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  718=>x"6600",	-- 0110011000000000  shr	r0, r0, 3
  719=>x"BBE8",	-- 1011101111101000  brieq	r5, put_sprite_16_aligned
  720=>x"062D",	-- 0000011000101101  dec	r5, r5
  721=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  722=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  723=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  724=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  725=>x"063F",	-- 0000011000111111  dec	r7, r7
  726=>x"D23B",	-- 1101001000111011  sw	r3, r7
  727=>x"0412",	-- 0000010000010010  inc	r2, r2
  728=>x"D011",	-- 1101000000010001  lw	r1, r2
  729=>x"CFF8",	-- 1100111111111000  li	r0, -1
  730=>x"3D40",	-- 0011110101000000  rsr	r0, r0, r5
  731=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  732=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  733=>x"D023",	-- 1101000000100011  lw	r3, r4
  734=>x"2600",	-- 0010011000000000  not	r0, r0
  735=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  736=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  737=>x"E421",	-- 1110010000100001  exw	r1, r4
  738=>x"0424",	-- 0000010000100100  inc	r4, r4
  739=>x"D011",	-- 1101000000010001  lw	r1, r2
  740=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  741=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  742=>x"D023",	-- 1101000000100011  lw	r3, r4
  743=>x"2600",	-- 0010011000000000  not	r0, r0
  744=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  745=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  746=>x"E421",	-- 1110010000100001  exw	r1, r4
  747=>x"0412",	-- 0000010000010010  inc	r2, r2
  748=>x"C098",	-- 1100000010011000  li	r0, 19
  749=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  750=>x"D03B",	-- 1101000000111011  lw	r3, r7
  751=>x"043F",	-- 0000010000111111  inc	r7, r7
  752=>x"061B",	-- 0000011000011011  dec	r3, r3
  753=>x"B91C",	-- 1011100100011100  brine	r3, put_sprite_16.loop
  754=>x"C005",	-- 1100000000000101  li	r5, 0
  755=>x"E383",	-- 1110001110000011  ba	-, r6
  756=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  757=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  758=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  759=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  760=>x"C005",	-- 1100000000000101  li	r5, 0
  761=>x"D020",	-- 1101000000100000  lw	r0, r4
  762=>x"D011",	-- 1101000000010001  lw	r1, r2
  763=>x"0412",	-- 0000010000010010  inc	r2, r2
  764=>x"2040",	-- 0010000001000000  and	r0, r0, r1
  765=>x"D011",	-- 1101000000010001  lw	r1, r2
  766=>x"0412",	-- 0000010000010010  inc	r2, r2
  767=>x"2240",	-- 0010001001000000  or	r0, r0, r1
  768=>x"E420",	-- 1110010000100000  exw	r0, r4
  769=>x"2040",	-- 0010000001000000  and	r0, r0, r1
  770=>x"222D",	-- 0010001000101101  or	r5, r5, r0
  771=>x"C0A0",	-- 1100000010100000  li	r0, 20
  772=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  773=>x"061B",	-- 0000011000011011  dec	r3, r3
  774=>x"AF5C",	-- 1010111101011100  brine	r3, put_sprite_16_aligned.loop
  775=>x"E383",	-- 1110001110000011  ba	-, r6
  776=>x"C07D",	-- 1100000001111101  li	r5, 15
  777=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  778=>x"6600",	-- 0110011000000000  shr	r0, r0, 3
  779=>x"BA68",	-- 1011101001101000  brieq	r5, put_sprite_16_masked_aligned
  780=>x"062D",	-- 0000011000101101  dec	r5, r5
  781=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  782=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  783=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  784=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  785=>x"063F",	-- 0000011000111111  dec	r7, r7
  786=>x"D23E",	-- 1101001000111110  sw	r6, r7
  787=>x"102E",	-- 0001000000101110  mova	r6, r5
  788=>x"C005",	-- 1100000000000101  li	r5, 0
  789=>x"063F",	-- 0000011000111111  dec	r7, r7
  790=>x"D23B",	-- 1101001000111011  sw	r3, r7
  791=>x"063F",	-- 0000011000111111  dec	r7, r7
  792=>x"D23B",	-- 1101001000111011  sw	r3, r7
  793=>x"D010",	-- 1101000000010000  lw	r0, r2
  794=>x"3980",	-- 0011100110000000  rrr	r0, r0, r6
  795=>x"0412",	-- 0000010000010010  inc	r2, r2
  796=>x"D011",	-- 1101000000010001  lw	r1, r2
  797=>x"3989",	-- 0011100110001001  rrr	r1, r1, r6
  798=>x"CFFD",	-- 1100111111111101  li	r5, -1
  799=>x"3DAD",	-- 0011110110101101  rsr	r5, r5, r6
  800=>x"2149",	-- 0010000101001001  and	r1, r1, r5
  801=>x"D023",	-- 1101000000100011  lw	r3, r4
  802=>x"262D",	-- 0010011000101101  not	r5, r5
  803=>x"222D",	-- 0010001000101101  or	r5, r5, r0
  804=>x"215B",	-- 0010000101011011  and	r3, r3, r5
  805=>x"225B",	-- 0010001001011011  or	r3, r3, r1
  806=>x"E423",	-- 1110010000100011  exw	r3, r4
  807=>x"205B",	-- 0010000001011011  and	r3, r3, r1
  808=>x"D03D",	-- 1101000000111101  lw	r5, r7
  809=>x"043F",	-- 0000010000111111  inc	r7, r7
  810=>x"22ED",	-- 0010001011101101  or	r5, r5, r3
  811=>x"0424",	-- 0000010000100100  inc	r4, r4
  812=>x"063F",	-- 0000011000111111  dec	r7, r7
  813=>x"D23B",	-- 1101001000111011  sw	r3, r7
  814=>x"D011",	-- 1101000000010001  lw	r1, r2
  815=>x"3989",	-- 0011100110001001  rrr	r1, r1, r6
  816=>x"CFFD",	-- 1100111111111101  li	r5, -1
  817=>x"3DAD",	-- 0011110110101101  rsr	r5, r5, r6
  818=>x"262D",	-- 0010011000101101  not	r5, r5
  819=>x"2149",	-- 0010000101001001  and	r1, r1, r5
  820=>x"D023",	-- 1101000000100011  lw	r3, r4
  821=>x"262D",	-- 0010011000101101  not	r5, r5
  822=>x"222D",	-- 0010001000101101  or	r5, r5, r0
  823=>x"215B",	-- 0010000101011011  and	r3, r3, r5
  824=>x"225B",	-- 0010001001011011  or	r3, r3, r1
  825=>x"E423",	-- 1110010000100011  exw	r3, r4
  826=>x"205B",	-- 0010000001011011  and	r3, r3, r1
  827=>x"D03D",	-- 1101000000111101  lw	r5, r7
  828=>x"043F",	-- 0000010000111111  inc	r7, r7
  829=>x"22ED",	-- 0010001011101101  or	r5, r5, r3
  830=>x"0412",	-- 0000010000010010  inc	r2, r2
  831=>x"C098",	-- 1100000010011000  li	r0, 19
  832=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  833=>x"D03B",	-- 1101000000111011  lw	r3, r7
  834=>x"043F",	-- 0000010000111111  inc	r7, r7
  835=>x"061B",	-- 0000011000011011  dec	r3, r3
  836=>x"B45C",	-- 1011010001011100  brine	r3, put_sprite_16_masked.loop
  837=>x"D03E",	-- 1101000000111110  lw	r6, r7
  838=>x"043F",	-- 0000010000111111  inc	r7, r7
  839=>x"E383",	-- 1110001110000011  ba	-, r6
  840=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  841=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  842=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  843=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  844=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  845=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  846=>x"C0A5",	-- 1100000010100101  li	r5, 20
  847=>x"8404",	-- 1000010000000100  brine	r0, put_sprite_8_aligned.loop1
  848=>x"D010",	-- 1101000000010000  lw	r0, r2
  849=>x"D021",	-- 1101000000100001  lw	r1, r4
  850=>x"1A41",	-- 0001101001000001  mixhl	r1, r0, r1
  851=>x"D221",	-- 1101001000100001  sw	r1, r4
  852=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  853=>x"061B",	-- 0000011000011011  dec	r3, r3
  854=>x"E398",	-- 1110001110011000  baeq	r3, r6
  855=>x"D021",	-- 1101000000100001  lw	r1, r4
  856=>x"1E41",	-- 0001111001000001  mixll	r1, r0, r1
  857=>x"D221",	-- 1101001000100001  sw	r1, r4
  858=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  859=>x"0412",	-- 0000010000010010  inc	r2, r2
  860=>x"061B",	-- 0000011000011011  dec	r3, r3
  861=>x"E398",	-- 1110001110011000  baeq	r3, r6
  862=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop0
  863=>x"D010",	-- 1101000000010000  lw	r0, r2
  864=>x"D021",	-- 1101000000100001  lw	r1, r4
  865=>x"1809",	-- 0001100000001001  mixhh	r1, r1, r0
  866=>x"D221",	-- 1101001000100001  sw	r1, r4
  867=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  868=>x"061B",	-- 0000011000011011  dec	r3, r3
  869=>x"E398",	-- 1110001110011000  baeq	r3, r6
  870=>x"D021",	-- 1101000000100001  lw	r1, r4
  871=>x"1A09",	-- 0001101000001001  mixhl	r1, r1, r0
  872=>x"D221",	-- 1101001000100001  sw	r1, r4
  873=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  874=>x"0412",	-- 0000010000010010  inc	r2, r2
  875=>x"061B",	-- 0000011000011011  dec	r3, r3
  876=>x"E398",	-- 1110001110011000  baeq	r3, r6
  877=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop1
  878=>x"C03D",	-- 1100000000111101  li	r5, 7
  879=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  880=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  881=>x"B5E8",	-- 1011010111101000  brieq	r5, put_sprite_8_aligned
  882=>x"062D",	-- 0000011000101101  dec	r5, r5
  883=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  884=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  885=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  886=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  887=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  888=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  889=>x"8A04",	-- 1000101000000100  brine	r0, put_sprite_8.loop1
  890=>x"D010",	-- 1101000000010000  lw	r0, r2
  891=>x"063F",	-- 0000011000111111  dec	r7, r7
  892=>x"D23A",	-- 1101001000111010  sw	r2, r7
  893=>x"C802",	-- 1100100000000010  li	r2, 0x100
  894=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  895=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  896=>x"D021",	-- 1101000000100001  lw	r1, r4
  897=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  898=>x"2612",	-- 0010011000010010  not	r2, r2
  899=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  900=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  901=>x"D221",	-- 1101001000100001  sw	r1, r4
  902=>x"C0A1",	-- 1100000010100001  li	r1, 20
  903=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  904=>x"D03A",	-- 1101000000111010  lw	r2, r7
  905=>x"043F",	-- 0000010000111111  inc	r7, r7
  906=>x"061B",	-- 0000011000011011  dec	r3, r3
  907=>x"E398",	-- 1110001110011000  baeq	r3, r6
  908=>x"D010",	-- 1101000000010000  lw	r0, r2
  909=>x"063F",	-- 0000011000111111  dec	r7, r7
  910=>x"D23A",	-- 1101001000111010  sw	r2, r7
  911=>x"1E00",	-- 0001111000000000  mixll	r0, r0, r0
  912=>x"C802",	-- 1100100000000010  li	r2, 0x100
  913=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  914=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  915=>x"D021",	-- 1101000000100001  lw	r1, r4
  916=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  917=>x"2612",	-- 0010011000010010  not	r2, r2
  918=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  919=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  920=>x"D221",	-- 1101001000100001  sw	r1, r4
  921=>x"C0A1",	-- 1100000010100001  li	r1, 20
  922=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  923=>x"D03A",	-- 1101000000111010  lw	r2, r7
  924=>x"043F",	-- 0000010000111111  inc	r7, r7
  925=>x"0412",	-- 0000010000010010  inc	r2, r2
  926=>x"061B",	-- 0000011000011011  dec	r3, r3
  927=>x"E398",	-- 1110001110011000  baeq	r3, r6
  928=>x"B683",	-- 1011011010000011  bri	-, put_sprite_8.loop0
  929=>x"D010",	-- 1101000000010000  lw	r0, r2
  930=>x"063F",	-- 0000011000111111  dec	r7, r7
  931=>x"D23A",	-- 1101001000111010  sw	r2, r7
  932=>x"063F",	-- 0000011000111111  dec	r7, r7
  933=>x"D23B",	-- 1101001000111011  sw	r3, r7
  934=>x"C802",	-- 1100100000000010  li	r2, 0x100
  935=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  936=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  937=>x"2080",	-- 0010000010000000  and	r0, r0, r2
  938=>x"D021",	-- 1101000000100001  lw	r1, r4
  939=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
  940=>x"261B",	-- 0010011000011011  not	r3, r3
  941=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  942=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
  943=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  944=>x"D221",	-- 1101001000100001  sw	r1, r4
  945=>x"0424",	-- 0000010000100100  inc	r4, r4
  946=>x"D021",	-- 1101000000100001  lw	r1, r4
  947=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  948=>x"261B",	-- 0010011000011011  not	r3, r3
  949=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  950=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
  951=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  952=>x"D221",	-- 1101001000100001  sw	r1, r4
  953=>x"C099",	-- 1100000010011001  li	r1, 19
  954=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  955=>x"D03B",	-- 1101000000111011  lw	r3, r7
  956=>x"043F",	-- 0000010000111111  inc	r7, r7
  957=>x"D03A",	-- 1101000000111010  lw	r2, r7
  958=>x"043F",	-- 0000010000111111  inc	r7, r7
  959=>x"061B",	-- 0000011000011011  dec	r3, r3
  960=>x"E398",	-- 1110001110011000  baeq	r3, r6
  961=>x"D010",	-- 1101000000010000  lw	r0, r2
  962=>x"4E00",	-- 0100111000000000  shl	r0, r0, 7
  963=>x"063F",	-- 0000011000111111  dec	r7, r7
  964=>x"D23A",	-- 1101001000111010  sw	r2, r7
  965=>x"063F",	-- 0000011000111111  dec	r7, r7
  966=>x"D23B",	-- 1101001000111011  sw	r3, r7
  967=>x"C802",	-- 1100100000000010  li	r2, 0x100
  968=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  969=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  970=>x"2080",	-- 0010000010000000  and	r0, r0, r2
  971=>x"D021",	-- 1101000000100001  lw	r1, r4
  972=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
  973=>x"261B",	-- 0010011000011011  not	r3, r3
  974=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  975=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
  976=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  977=>x"D221",	-- 1101001000100001  sw	r1, r4
  978=>x"0424",	-- 0000010000100100  inc	r4, r4
  979=>x"D021",	-- 1101000000100001  lw	r1, r4
  980=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  981=>x"261B",	-- 0010011000011011  not	r3, r3
  982=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  983=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
  984=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  985=>x"D221",	-- 1101001000100001  sw	r1, r4
  986=>x"C099",	-- 1100000010011001  li	r1, 19
  987=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  988=>x"D03B",	-- 1101000000111011  lw	r3, r7
  989=>x"043F",	-- 0000010000111111  inc	r7, r7
  990=>x"D03A",	-- 1101000000111010  lw	r2, r7
  991=>x"043F",	-- 0000010000111111  inc	r7, r7
  992=>x"0412",	-- 0000010000010010  inc	r2, r2
  993=>x"061B",	-- 0000011000011011  dec	r3, r3
  994=>x"E398",	-- 1110001110011000  baeq	r3, r6
  995=>x"AF83",	-- 1010111110000011  bri	-, put_sprite_8.loop1
    others => x"0000"
    );
begin
  process(CLK)
  begin
    if (CLK'event AND CLK='1') then
      D <= m(to_integer(unsigned(AD)));
    end if;
  end process;
end Behavioral;
