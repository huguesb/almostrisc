----------------------------------------------------------------------------------
--
-- File retrieved, on 07/02/2010, from :
-- http://sebastien-viardot.imag.fr/Enseignements/Archi1A2s/sources/ROMPROG.vhd
--
-- Slightly altered to get rid of vendor-specific packages and adjust formatting
-- Now auto-filled by asrom script
--
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROMPROG is
  Port ( AD : in  STD_LOGIC_VECTOR (12 downto 0);
         D : out  STD_LOGIC_VECTOR (15 downto 0);
         CLK : in STD_LOGIC);
end ROMPROG;

architecture Behavioral of ROMPROG is
  constant low_address: natural := 0;
  constant high_address: natural := 8192;
  subtype octet is std_logic_vector( 15 downto 0 );
  type zone_memoire is
    array (natural range low_address to high_address-1) of octet;
  constant m: zone_memoire:= (
    0=>x"FFF7",	-- 1111111111110111  liw	r7, IRQ_mask
    1=>x"2000",	-- 0010000000000000  
    2=>x"F8C0",	-- 1111100011000000  bai	-, os_init
    3=>x"0100",	-- 0000000100000000  
   16=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_ack
   17=>x"2002",	-- 0010000000000010  
   18=>x"D001",	-- 1101000000000001  lw	r1, r0
   19=>x"F54A",	-- 1111010101001010  bspl	r2, r1, 5
   20=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_error
   21=>x"0050",	-- 0000000001010000  
   22=>x"F4CA",	-- 1111010011001010  bspl	r2, r1, 3
   23=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_kbd
   24=>x"0060",	-- 0000000001100000  
   25=>x"F40A",	-- 1111010000001010  bspl	r2, r1, 0
   26=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_tmr
   27=>x"0040",	-- 0000000001000000  
   28=>x"D201",	-- 1101001000000001  sw	r1, r0
   29=>x"FFFE",	-- 1111111111111110  reti
   64=>x"263F",	-- 0010011000111111  not r7, r7
   65=>x"D7C0",	-- 1101011111000000  out	r7
   66=>x"E383",	-- 1110001110000011  ba	-, r6
   80=>x"25FF",	-- 0010010111111111  xor	r7, r7, r7
   81=>x"D7C0",	-- 1101011111000000  out	r7
   82=>x"E383",	-- 1110001110000011  ba	-, r6
   96=>x"FFF2",	-- 1111111111110010  liw	r2, PS2_rx
   97=>x"2004",	-- 0010000000000100  
   98=>x"D012",	-- 1101000000010010  lw	r2, r2
   99=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map + 8
  100=>x"1808",	-- 0001100000001000  
  101=>x"D01B",	-- 1101000000011011  lw	r3, r3
  102=>x"1EBF",	-- 0001111010111111  mixll	r7, r7, r2
  103=>x"C784",	-- 1100011110000100  li	r4, 0xF0
  104=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  105=>x"8B20",	-- 1000101100100000  brieq	r4, int_kbd.release
  106=>x"C704",	-- 1100011100000100  li	r4, 0xE0
  107=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  108=>x"88E0",	-- 1000100011100000  brieq	r4, int_kbd.extended
  109=>x"FFF5",	-- 1111111111110101  liw	r5, paper_keys - 1
  110=>x"16BF",	-- 0001011010111111  
  111=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  112=>x"80E0",	-- 1000000011100000  brieq	r4, $+3
  113=>x"FFF5",	-- 1111111111110101  liw	r5, paper_keys + 11 - 1
  114=>x"16CA",	-- 0001011011001010  
  115=>x"042D",	-- 0000010000101101  inc	r5, r5
  116=>x"D02C",	-- 1101000000101100  lw	r4, r5
  117=>x"8560",	-- 1000010101100000  brieq	r4, scan_code_mismatch
  118=>x"6E24",	-- 0110111000100100  shr	r4, r4, 7
  119=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  120=>x"BEE4",	-- 1011111011100100  brine	r4, scan_code_loop
  121=>x"D02A",	-- 1101000000101010  lw	r2, r5
  122=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  123=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  124=>x"741B",	-- 0111010000011011  shr	r3, r3, 10
  125=>x"C00D",	-- 1100000000001101  li	r5, 1
  126=>x"0612",	-- 0000011000010010  dec	r2, r2
  127=>x"3AAA",	-- 0011101010101010  rrl	r2, r5, r2
  128=>x"FFF5",	-- 1111111111110101  liw	r5, key_press_map
  129=>x"1800",	-- 0001100000000000  
  130=>x"08ED",	-- 0000100011101101  add	r5, r5, r3
  131=>x"D02B",	-- 1101000000101011  lw	r3, r5
  132=>x"80E4",	-- 1000000011100100  brine	r4, scan_code_release
  133=>x"229B",	-- 0010001010011011  or	r3, r3, r2
  134=>x"80C3",	-- 1000000011000011  bri	-, scan_code_notify
  135=>x"2612",	-- 0010011000010010  not	r2, r2
  136=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  137=>x"D22B",	-- 1101001000101011  sw	r3, r5
  138=>x"C003",	-- 1100000000000011  li	r3, 0
  139=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  140=>x"1808",	-- 0001100000001000  
  141=>x"D223",	-- 1101001000100011  sw	r3, r4
  142=>x"E383",	-- 1110001110000011  ba	-, r6
  143=>x"C014",	-- 1100000000010100  li	r4, 2
  144=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  145=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  146=>x"1808",	-- 0001100000001000  
  147=>x"D223",	-- 1101001000100011  sw	r3, r4
  148=>x"E383",	-- 1110001110000011  ba	-, r6
  149=>x"C00C",	-- 1100000000001100  li	r4, 1
  150=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  151=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  152=>x"1808",	-- 0001100000001000  
  153=>x"D223",	-- 1101001000100011  sw	r3, r4
  154=>x"E383",	-- 1110001110000011  ba	-, r6
  256=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_mask
  257=>x"2000",	-- 0010000000000000  
  258=>x"C0C9",	-- 1100000011001001  li	r1, 0x19
  259=>x"D201",	-- 1101001000000001  sw	r1, r0
  260=>x"0400",	-- 0000010000000000  inc	r0, r0
  261=>x"CFF9",	-- 1100111111111001  li	r1, -1
  262=>x"D201",	-- 1101001000000001  sw	r1, r0
  263=>x"C03A",	-- 1100000000111010  li	r2, 7
  264=>x"0880",	-- 0000100010000000  add	r0, r0, r2
  265=>x"C0EA",	-- 1100000011101010  li	r2, 0x1D
  266=>x"D202",	-- 1101001000000010  sw	r2, r0
  267=>x"0400",	-- 0000010000000000  inc	r0, r0
  268=>x"C07A",	-- 1100000001111010  li	r2, 15
  269=>x"D202",	-- 1101001000000010  sw	r2, r0
  270=>x"FFF0",	-- 1111111111110000  liw	r0, key_press_map
  271=>x"1800",	-- 0001100000000000  
  272=>x"C001",	-- 1100000000000001  li	r1, 0
  273=>x"C042",	-- 1100000001000010  li	r2, 8
  274=>x"D201",	-- 1101001000000001  sw	r1, r0
  275=>x"0400",	-- 0000010000000000  inc	r0, r0
  276=>x"0612",	-- 0000011000010010  dec	r2, r2
  277=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  278=>x"C0F3",	-- 1100000011110011  li	r3, 30
  279=>x"CFFA",	-- 1100111111111010  li	r2, -1
  280=>x"D21A",	-- 1101001000011010  sw	r2, r3
  281=>x"8083",	-- 1000000010000011  bri	-, PaperGameStart
  282=>x"8003",	-- 1000000000000011  bri	-, PaperMenuLoop
  283=>x"FFF0",	-- 1111111111110000  liw	r0, paper_dir
  284=>x"173C",	-- 0001011100111100  
  285=>x"C001",	-- 1100000000000001  li	r1, 0
  286=>x"D201",	-- 1101001000000001  sw	r1, r0
  287=>x"0400",	-- 0000010000000000  inc	r0, r0
  288=>x"FFF1",	-- 1111111111110001  liw	r1, 152 * 8
  289=>x"04C0",	-- 0000010011000000  
  290=>x"D201",	-- 1101001000000001  sw	r1, r0
  291=>x"0400",	-- 0000010000000000  inc	r0, r0
  292=>x"C001",	-- 1100000000000001  li	r1, 0
  293=>x"D201",	-- 1101001000000001  sw	r1, r0
  294=>x"0400",	-- 0000010000000000  inc	r0, r0
  295=>x"FFF1",	-- 1111111111110001  liw	r1, 128 * 8
  296=>x"0400",	-- 0000010000000000  
  297=>x"D201",	-- 1101001000000001  sw	r1, r0
  298=>x"0400",	-- 0000010000000000  inc	r0, r0
  299=>x"C001",	-- 1100000000000001  li	r1, 0
  300=>x"D201",	-- 1101001000000001  sw	r1, r0
  301=>x"0400",	-- 0000010000000000  inc	r0, r0
  302=>x"C029",	-- 1100000000101001  li	r1, 5
  303=>x"D201",	-- 1101001000000001  sw	r1, r0
  304=>x"0400",	-- 0000010000000000  inc	r0, r0
  305=>x"C011",	-- 1100000000010001  li	r1, 2
  306=>x"D201",	-- 1101001000000001  sw	r1, r0
  307=>x"0400",	-- 0000010000000000  inc	r0, r0
  308=>x"C000",	-- 1100000000000000  li	r0, 0
  309=>x"CFF9",	-- 1100111111111001  li	r1, -1
  310=>x"C0A2",	-- 1100000010100010  li	r2, 20
  311=>x"D201",	-- 1101001000000001  sw	r1, r0
  312=>x"0400",	-- 0000010000000000  inc	r0, r0
  313=>x"0612",	-- 0000011000010010  dec	r2, r2
  314=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  315=>x"C001",	-- 1100000000000001  li	r1, 0
  316=>x"FFF2",	-- 1111111111110010  liw	r2, 18*20
  317=>x"0168",	-- 0000000101101000  
  318=>x"D201",	-- 1101001000000001  sw	r1, r0
  319=>x"0400",	-- 0000010000000000  inc	r0, r0
  320=>x"0612",	-- 0000011000010010  dec	r2, r2
  321=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  322=>x"CFF9",	-- 1100111111111001  li	r1, -1
  323=>x"C0A2",	-- 1100000010100010  li	r2, 20
  324=>x"D201",	-- 1101001000000001  sw	r1, r0
  325=>x"0400",	-- 0000010000000000  inc	r0, r0
  326=>x"0612",	-- 0000011000010010  dec	r2, r2
  327=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  328=>x"C020",	-- 1100000000100000  li	r0, 4
  329=>x"C029",	-- 1100000000101001  li	r1, 5
  330=>x"FFF2",	-- 1111111111110010  liw	r2, paper_title
  331=>x"1744",	-- 0001011101000100  
  332=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  333=>x"024A",	-- 0000001001001010  
  334=>x"C778",	-- 1100011101111000  li	r0, 239
  335=>x"C009",	-- 1100000000001001  li	r1, 1
  336=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud
  337=>x"1720",	-- 0001011100100000  
  338=>x"C043",	-- 1100000001000011  li	r3, 8
  339=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  340=>x"02F4",	-- 0000001011110100  
  341=>x"C0F8",	-- 1100000011111000  li	r0, 31
  342=>x"C009",	-- 1100000000001001  li	r1, 1
  343=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed + 1
  344=>x"1741",	-- 0001011101000001  
  345=>x"D012",	-- 1101000000010010  lw	r2, r2
  346=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum
  347=>x"0279",	-- 0000001001111001  
  348=>x"C120",	-- 1100000100100000  li	r0, 36
  349=>x"C009",	-- 1100000000001001  li	r1, 1
  350=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  351=>x"174A",	-- 0001011101001010  
  352=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  353=>x"024A",	-- 0000001001001010  
  354=>x"C778",	-- 1100011101111000  li	r0, 239
  355=>x"C051",	-- 1100000001010001  li	r1, 10
  356=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud + 4
  357=>x"1724",	-- 0001011100100100  
  358=>x"C043",	-- 1100000001000011  li	r3, 8
  359=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  360=>x"02F4",	-- 0000001011110100  
  361=>x"C0F8",	-- 1100000011111000  li	r0, 31
  362=>x"C051",	-- 1100000001010001  li	r1, 10
  363=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed + 2
  364=>x"1742",	-- 0001011101000010  
  365=>x"D012",	-- 1101000000010010  lw	r2, r2
  366=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum
  367=>x"0279",	-- 0000001001111001  
  368=>x"C120",	-- 1100000100100000  li	r0, 36
  369=>x"C051",	-- 1100000001010001  li	r1, 10
  370=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  371=>x"174A",	-- 0001011101001010  
  372=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  373=>x"024A",	-- 0000001001001010  
  374=>x"FFF0",	-- 1111111111110000  liw	r0, 20*20
  375=>x"0190",	-- 0000000110010000  
  376=>x"C001",	-- 1100000000000001  li	r1, 0
  377=>x"FFF2",	-- 1111111111110010  liw	r2, 220*20
  378=>x"1130",	-- 0001000100110000  
  379=>x"D201",	-- 1101001000000001  sw	r1, r0
  380=>x"0400",	-- 0000010000000000  inc	r0, r0
  381=>x"0612",	-- 0000011000010010  dec	r2, r2
  382=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  383=>x"FFF5",	-- 1111111111110101  liw	r5, paper_tilemap
  384=>x"1780",	-- 0001011110000000  
  385=>x"D02C",	-- 1101000000101100  lw	r4, r5
  386=>x"042D",	-- 0000010000101101  inc	r5, r5
  387=>x"8720",	-- 1000011100100000  brieq	r4, PaperGameTileSkip
  388=>x"063F",	-- 0000011000111111  dec	r7, r7
  389=>x"D23D",	-- 1101001000111101  sw	r5, r7
  390=>x"FFF3",	-- 1111111111110011  liw	r3, paper_tilemap
  391=>x"1780",	-- 0001011110000000  
  392=>x"0AEB",	-- 0000101011101011  sub	r3, r5, r3
  393=>x"6E20",	-- 0110111000100000  shr	r0, r4, 7
  394=>x"6219",	-- 0110001000011001  shr	r1, r3, 1
  395=>x"4409",	-- 0100010000001001  shl	r1, r1, 2
  396=>x"FFF2",	-- 1111111111110010  liw	r2, paper_pos + 1
  397=>x"173E",	-- 0001011100111110  
  398=>x"D012",	-- 1101000000010010  lw	r2, r2
  399=>x"6412",	-- 0110010000010010  shr	r2, r2, 2
  400=>x"C03B",	-- 1100000000111011  li	r3, 7
  401=>x"20D2",	-- 0010000011010010  and	r2, r2, r3
  402=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  403=>x"4E24",	-- 0100111000100100  shl	r4, r4, 7
  404=>x"6E24",	-- 0110111000100100  shr	r4, r4, 7
  405=>x"C00B",	-- 1100000000001011  li	r3, 1
  406=>x"FB06",	-- 1111101100000110  bailne	r0, r6, put_tile
  407=>x"01F6",	-- 0000000111110110  
  408=>x"C013",	-- 1100000000010011  li	r3, 2
  409=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_tile
  410=>x"01F6",	-- 0000000111110110  
  411=>x"0624",	-- 0000011000100100  dec	r4, r4
  412=>x"BF64",	-- 1011111101100100  brine	r4, PaperGameSegmentLoop
  413=>x"D03D",	-- 1101000000111101  lw	r5, r7
  414=>x"043F",	-- 0000010000111111  inc	r7, r7
  415=>x"FFF4",	-- 1111111111110100  liw r4, paper_tilemap + 125
  416=>x"17FD",	-- 0001011111111101  
  417=>x"0B2C",	-- 0000101100101100  sub	r4, r5, r4
  418=>x"B7E5",	-- 1011011111100101  brilt	r4, PaperGameTileLoop
  419=>x"FFF3",	-- 1111111111110011  liw	r3, paper_speed
  420=>x"1740",	-- 0001011101000000  
  421=>x"D01C",	-- 1101000000011100  lw	r4, r3
  422=>x"F7E5",	-- 1111011111100101  bspl	r5, r4, 15
  423=>x"2564",	-- 0010010101100100  xor	r4, r4, r5
  424=>x"6424",	-- 0110010000100100  shr	r4, r4, 2
  425=>x"2564",	-- 0010010101100100  xor	r4, r4, r5
  426=>x"FFF3",	-- 1111111111110011  liw	r3, paper_pos
  427=>x"173D",	-- 0001011100111101  
  428=>x"D018",	-- 1101000000011000  lw	r0, r3
  429=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  430=>x"FFF2",	-- 1111111111110010  liw	r2, paper_sprites
  431=>x"16F0",	-- 0001011011110000  
  432=>x"4624",	-- 0100011000100100  shl	r4, r4, 3
  433=>x"0912",	-- 0000100100010010  add	r2, r2, r4
  434=>x"C161",	-- 1100000101100001  li	r1, 44
  435=>x"C083",	-- 1100000010000011  li	r3, 16
  436=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_16
  437=>x"02A8",	-- 0000001010101000  
  438=>x"C028",	-- 1100000000101000  li	r0, 5
  439=>x"C001",	-- 1100000000000001  li	r1, 0
  440=>x"8043",	-- 1000000001000011  bri	-, $+1
  441=>x"8043",	-- 1000000001000011  bri	-, $+1
  442=>x"0609",	-- 0000011000001001  dec	r1, r1
  443=>x"BF4C",	-- 1011111101001100  brine	r1, $-3
  444=>x"0600",	-- 0000011000000000  dec	r0, r0
  445=>x"BE84",	-- 1011111010000100  brine	r0, $-6
  446=>x"FFF2",	-- 1111111111110010  liw	r2, paper_pos
  447=>x"173D",	-- 0001011100111101  
  448=>x"FFF3",	-- 1111111111110011  liw	r3, paper_speed
  449=>x"1740",	-- 0001011101000000  
  450=>x"D010",	-- 1101000000010000  lw	r0, r2
  451=>x"D019",	-- 1101000000011001  lw	r1, r3
  452=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  453=>x"D210",	-- 1101001000010000  sw	r0, r2
  454=>x"0412",	-- 0000010000010010  inc	r2, r2
  455=>x"041B",	-- 0000010000011011  inc	r3, r3
  456=>x"D010",	-- 1101000000010000  lw	r0, r2
  457=>x"D019",	-- 1101000000011001  lw	r1, r3
  458=>x"C1FC",	-- 1100000111111100  li	r4, 0x3F
  459=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  460=>x"2101",	-- 0010000100000001  and	r1, r0, r4
  461=>x"2624",	-- 0010011000100100  not	r4, r4
  462=>x"2100",	-- 0010000100000000  and	r0, r0, r4
  463=>x"D211",	-- 1101001000010001  sw	r1, r2
  464=>x"8300",	-- 1000001100000000  brieq	r0, PaperGameSkipScroll
  465=>x"FFF0",	-- 1111111111110000  liw	r0, paper_tilemap
  466=>x"1780",	-- 0001011110000000  
  467=>x"C021",	-- 1100000000100001  li	r1, 4
  468=>x"0841",	-- 0000100001000001  add	r1, r0, r1
  469=>x"C302",	-- 1100001100000010  li	r2, 24*4
  470=>x"D00B",	-- 1101000000001011  lw	r3, r1
  471=>x"D203",	-- 1101001000000011  sw	r3, r0
  472=>x"0400",	-- 0000010000000000  inc	r0, r0
  473=>x"0409",	-- 0000010000001001  inc	r1, r1
  474=>x"0612",	-- 0000011000010010  dec	r2, r2
  475=>x"BED4",	-- 1011111011010100  brine	r2, PaperGameScrollLoop
  476=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  477=>x"1800",	-- 0001100000000000  
  478=>x"D01B",	-- 1101000000011011  lw	r3, r3
  479=>x"A5D8",	-- 1010010111011000  brieq	r3, PaperGameRedrawContent
  480=>x"F7DC",	-- 1111011111011100  bspl	r4, r3, 15
  481=>x"8524",	-- 1000010100100100  brine	r4, PaperGameQuit
  482=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  483=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveUp
  484=>x"F49C",	-- 1111010010011100  bspl	r4, r3, 2
  485=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveDOWN
  486=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  487=>x"81A0",	-- 1000000110100000  brieq	r4, PaperNoMoveLEFT
  488=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  489=>x"1740",	-- 0001011101000000  
  490=>x"D010",	-- 1101000000010000  lw	r0, r2
  491=>x"0600",	-- 0000011000000000  dec	r0, r0
  492=>x"D210",	-- 1101001000010000  sw	r0, r2
  493=>x"F4DC",	-- 1111010011011100  bspl	r4, r3, 3
  494=>x"81A0",	-- 1000000110100000  brieq	r4, PaperNoMoveRIGHT
  495=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  496=>x"1740",	-- 0001011101000000  
  497=>x"D010",	-- 1101000000010000  lw	r0, r2
  498=>x"0400",	-- 0000010000000000  inc	r0, r0
  499=>x"D210",	-- 1101001000010000  sw	r0, r2
  500=>x"A083",	-- 1010000010000011  bri	-, PaperGameRedrawContent
  501=>x"FFFF",	-- 1111111111111111  reset
  502=>x"063F",	-- 0000011000111111  dec	r7, r7
  503=>x"D238",	-- 1101001000111000  sw	r0, r7
  504=>x"063F",	-- 0000011000111111  dec	r7, r7
  505=>x"D239",	-- 1101001000111001  sw	r1, r7
  506=>x"063F",	-- 0000011000111111  dec	r7, r7
  507=>x"D23A",	-- 1101001000111010  sw	r2, r7
  508=>x"063F",	-- 0000011000111111  dec	r7, r7
  509=>x"D23B",	-- 1101001000111011  sw	r3, r7
  510=>x"063F",	-- 0000011000111111  dec	r7, r7
  511=>x"D23C",	-- 1101001000111100  sw	r4, r7
  512=>x"063F",	-- 0000011000111111  dec	r7, r7
  513=>x"D23D",	-- 1101001000111101  sw	r5, r7
  514=>x"063F",	-- 0000011000111111  dec	r7, r7
  515=>x"D23E",	-- 1101001000111110  sw	r6, r7
  516=>x"FFF2",	-- 1111111111110010  liw	r2, paper_tiles
  517=>x"1730",	-- 0001011100110000  
  518=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  519=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  520=>x"C043",	-- 1100000001000011  li	r3, 8
  521=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  522=>x"02CE",	-- 0000001011001110  
  523=>x"D03E",	-- 1101000000111110  lw	r6, r7
  524=>x"043F",	-- 0000010000111111  inc	r7, r7
  525=>x"D03D",	-- 1101000000111101  lw	r5, r7
  526=>x"043F",	-- 0000010000111111  inc	r7, r7
  527=>x"D03C",	-- 1101000000111100  lw	r4, r7
  528=>x"043F",	-- 0000010000111111  inc	r7, r7
  529=>x"D03B",	-- 1101000000111011  lw	r3, r7
  530=>x"043F",	-- 0000010000111111  inc	r7, r7
  531=>x"D03A",	-- 1101000000111010  lw	r2, r7
  532=>x"043F",	-- 0000010000111111  inc	r7, r7
  533=>x"D039",	-- 1101000000111001  lw	r1, r7
  534=>x"043F",	-- 0000010000111111  inc	r7, r7
  535=>x"D038",	-- 1101000000111000  lw	r0, r7
  536=>x"043F",	-- 0000010000111111  inc	r7, r7
  537=>x"0400",	-- 0000010000000000  inc	r0, r0
  538=>x"E383",	-- 1110001110000011  ba	-, r6
  539=>x"C750",	-- 1100011101010000  li	r0, 234
  540=>x"C1C2",	-- 1100000111000010  li	r2, 56
  541=>x"FAC6",	-- 1111101011000110  bail	-, r6, div_16_16
  542=>x"0233",	-- 0000001000110011  
  543=>x"C448",	-- 1100010001001000  li	r0, 137
  544=>x"C472",	-- 1100010001110010  li	r2, 142
  545=>x"FAC6",	-- 1111101011000110  bail	-, r6, mult_16_16
  546=>x"0227",	-- 0000001000100111  
  547=>x"C03A",	-- 1100000000111010  li r2, 7
  548=>x"FAC6",	-- 1111101011000110  bail	-, r6, fact_16
  549=>x"023E",	-- 0000001000111110  
  550=>x"FFFF",	-- 1111111111111111  reset
  551=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  552=>x"2524",	-- 0010010100100100  xor	r4, r4, r4
  553=>x"C085",	-- 1100000010000101  li	r5, 16
  554=>x"0849",	-- 0000100001001001  add	r1, r1, r1
  555=>x"0C00",	-- 0000110000000000  adc	r0, r0, r0
  556=>x"0EDB",	-- 0000111011011011  sbc	r3, r3, r3
  557=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  558=>x"08C9",	-- 0000100011001001  add	r1, r1, r3
  559=>x"0D00",	-- 0000110100000000  adc	r0, r0, r4
  560=>x"062D",	-- 0000011000101101  dec	r5, r5
  561=>x"BE6C",	-- 1011111001101100  brine	r5, mult_16_16.loop
  562=>x"E383",	-- 1110001110000011  ba	-, r6
  563=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  564=>x"C084",	-- 1100000010000100  li	r4, 16
  565=>x"0800",	-- 0000100000000000  add	r0, r0, r0
  566=>x"0C49",	-- 0000110001001001  adc	r1, r1, r1
  567=>x"0A8B",	-- 0000101010001011  sub	r3, r1, r2
  568=>x"80DD",	-- 1000000011011101  brilt	r3, div_16_16.skip
  569=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  570=>x"0400",	-- 0000010000000000  inc	r0, r0
  571=>x"0624",	-- 0000011000100100  dec	r4, r4
  572=>x"BE64",	-- 1011111001100100  brine	r4, div_16_16.loop
  573=>x"E383",	-- 1110001110000011  ba	-, r6
  574=>x"2400",	-- 0010010000000000  xor	r0, r0, r0
  575=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  576=>x"8250",	-- 1000001001010000  brieq	r2, fact_16.end
  577=>x"0409",	-- 0000010000001001  inc	r1, r1
  578=>x"1008",	-- 0001000000001000  mova	r0, r1
  579=>x"FAC6",	-- 1111101011000110  bail	-, r6, mult_16_16
  580=>x"0227",	-- 0000001000100111  
  581=>x"8104",	-- 1000000100000100  brine	r0, fact_16.overflow
  582=>x"0227",	-- 0000001000100111  
  583=>x"0612",	-- 0000011000010010  dec	r2, r2
  584=>x"BE94",	-- 1011111010010100  brine	r2, fact_16.loop
  585=>x"E383",	-- 1110001110000011  ba	-, r6
  586=>x"063F",	-- 0000011000111111  dec	r7, r7
  587=>x"D23E",	-- 1101001000111110  sw	r6, r7
  588=>x"D013",	-- 1101000000010011  lw	r3, r2
  589=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  590=>x"84D8",	-- 1000010011011000  brieq	r3, puts.end
  591=>x"063F",	-- 0000011000111111  dec	r7, r7
  592=>x"D23A",	-- 1101001000111010  sw	r2, r7
  593=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  594=>x"0264",	-- 0000001001100100  
  595=>x"D03A",	-- 1101000000111010  lw	r2, r7
  596=>x"043F",	-- 0000010000111111  inc	r7, r7
  597=>x"D013",	-- 1101000000010011  lw	r3, r2
  598=>x"4E1B",	-- 0100111000011011  shl	r3, r3, 7
  599=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  600=>x"8258",	-- 1000001001011000  brieq	r3, puts.end
  601=>x"063F",	-- 0000011000111111  dec	r7, r7
  602=>x"D23A",	-- 1101001000111010  sw	r2, r7
  603=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  604=>x"0264",	-- 0000001001100100  
  605=>x"D03A",	-- 1101000000111010  lw	r2, r7
  606=>x"043F",	-- 0000010000111111  inc	r7, r7
  607=>x"0412",	-- 0000010000010010  inc	r2, r2
  608=>x"BB03",	-- 1011101100000011  bri	-, puts.loop
  609=>x"D03E",	-- 1101000000111110  lw	r6, r7
  610=>x"043F",	-- 0000010000111111  inc	r7, r7
  611=>x"E383",	-- 1110001110000011  ba	-, r6
  612=>x"063F",	-- 0000011000111111  dec	r7, r7
  613=>x"D23E",	-- 1101001000111110  sw	r6, r7
  614=>x"063F",	-- 0000011000111111  dec	r7, r7
  615=>x"D238",	-- 1101001000111000  sw	r0, r7
  616=>x"063F",	-- 0000011000111111  dec	r7, r7
  617=>x"D239",	-- 1101001000111001  sw	r1, r7
  618=>x"FFF2",	-- 1111111111110010  liw	r2, font_map
  619=>x"12C0",	-- 0001001011000000  
  620=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  621=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  622=>x"C043",	-- 1100000001000011  li	r3, 8
  623=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  624=>x"02CE",	-- 0000001011001110  
  625=>x"D039",	-- 1101000000111001  lw	r1, r7
  626=>x"043F",	-- 0000010000111111  inc	r7, r7
  627=>x"D038",	-- 1101000000111000  lw	r0, r7
  628=>x"043F",	-- 0000010000111111  inc	r7, r7
  629=>x"0400",	-- 0000010000000000  inc	r0, r0
  630=>x"D03E",	-- 1101000000111110  lw	r6, r7
  631=>x"043F",	-- 0000010000111111  inc	r7, r7
  632=>x"E383",	-- 1110001110000011  ba	-, r6
  633=>x"063F",	-- 0000011000111111  dec	r7, r7
  634=>x"D23E",	-- 1101001000111110  sw	r6, r7
  635=>x"FFF4",	-- 1111111111110100  liw	r4, 10000
  636=>x"2710",	-- 0010011100010000  
  637=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  638=>x"028C",	-- 0000001010001100  
  639=>x"FFF4",	-- 1111111111110100  liw	r4, 1000
  640=>x"03E8",	-- 0000001111101000  
  641=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  642=>x"028C",	-- 0000001010001100  
  643=>x"C324",	-- 1100001100100100  li	r4, 100
  644=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  645=>x"028C",	-- 0000001010001100  
  646=>x"C054",	-- 1100000001010100  li	r4, 10
  647=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  648=>x"028C",	-- 0000001010001100  
  649=>x"D03E",	-- 1101000000111110  lw	r6, r7
  650=>x"043F",	-- 0000010000111111  inc	r7, r7
  651=>x"C00C",	-- 1100000000001100  li	r4, 1
  652=>x"C17B",	-- 1100000101111011  li	r3, 0x2F
  653=>x"041B",	-- 0000010000011011  inc	r3, r3
  654=>x"0B12",	-- 0000101100010010  sub	r2, r2, r4
  655=>x"BF91",	-- 1011111110010001  brige	r2, printnum.loop
  656=>x"0912",	-- 0000100100010010  add	r2, r2, r4
  657=>x"063F",	-- 0000011000111111  dec	r7, r7
  658=>x"D23E",	-- 1101001000111110  sw	r6, r7
  659=>x"063F",	-- 0000011000111111  dec	r7, r7
  660=>x"D23A",	-- 1101001000111010  sw	r2, r7
  661=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  662=>x"0264",	-- 0000001001100100  
  663=>x"D03A",	-- 1101000000111010  lw	r2, r7
  664=>x"043F",	-- 0000010000111111  inc	r7, r7
  665=>x"D03E",	-- 1101000000111110  lw	r6, r7
  666=>x"043F",	-- 0000010000111111  inc	r7, r7
  667=>x"E383",	-- 1110001110000011  ba	-, r6
  668=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  669=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  670=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  671=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  672=>x"C0A0",	-- 1100000010100000  li	r0, 20
  673=>x"D011",	-- 1101000000010001  lw	r1, r2
  674=>x"D221",	-- 1101001000100001  sw	r1, r4
  675=>x"0412",	-- 0000010000010010  inc	r2, r2
  676=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  677=>x"061B",	-- 0000011000011011  dec	r3, r3
  678=>x"BEDC",	-- 1011111011011100  brine	r3, put_sprite_16_aligned.loop
  679=>x"E383",	-- 1110001110000011  ba	-, r6
  680=>x"C07D",	-- 1100000001111101  li	r5, 15
  681=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  682=>x"6600",	-- 0110011000000000  shr	r0, r0, 3
  683=>x"BC68",	-- 1011110001101000  brieq	r5, put_sprite_16_aligned
  684=>x"062D",	-- 0000011000101101  dec	r5, r5
  685=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  686=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  687=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  688=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  689=>x"063F",	-- 0000011000111111  dec	r7, r7
  690=>x"D23B",	-- 1101001000111011  sw	r3, r7
  691=>x"D011",	-- 1101000000010001  lw	r1, r2
  692=>x"CFF8",	-- 1100111111111000  li	r0, -1
  693=>x"3D40",	-- 0011110101000000  rsr	r0, r0, r5
  694=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  695=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  696=>x"D023",	-- 1101000000100011  lw	r3, r4
  697=>x"2600",	-- 0010011000000000  not	r0, r0
  698=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  699=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  700=>x"D221",	-- 1101001000100001  sw	r1, r4
  701=>x"0424",	-- 0000010000100100  inc	r4, r4
  702=>x"D011",	-- 1101000000010001  lw	r1, r2
  703=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  704=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  705=>x"D023",	-- 1101000000100011  lw	r3, r4
  706=>x"2600",	-- 0010011000000000  not	r0, r0
  707=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  708=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  709=>x"D221",	-- 1101001000100001  sw	r1, r4
  710=>x"0412",	-- 0000010000010010  inc	r2, r2
  711=>x"C098",	-- 1100000010011000  li	r0, 19
  712=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  713=>x"D03B",	-- 1101000000111011  lw	r3, r7
  714=>x"043F",	-- 0000010000111111  inc	r7, r7
  715=>x"061B",	-- 0000011000011011  dec	r3, r3
  716=>x"B95C",	-- 1011100101011100  brine	r3, put_sprite_16.loop
  717=>x"E383",	-- 1110001110000011  ba	-, r6
  718=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  719=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  720=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  721=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  722=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  723=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  724=>x"C0A5",	-- 1100000010100101  li	r5, 20
  725=>x"8404",	-- 1000010000000100  brine	r0, put_sprite_8_aligned.loop1
  726=>x"D010",	-- 1101000000010000  lw	r0, r2
  727=>x"D021",	-- 1101000000100001  lw	r1, r4
  728=>x"1A41",	-- 0001101001000001  mixhl	r1, r0, r1
  729=>x"D221",	-- 1101001000100001  sw	r1, r4
  730=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  731=>x"061B",	-- 0000011000011011  dec	r3, r3
  732=>x"E398",	-- 1110001110011000  baeq	r3, r6
  733=>x"D021",	-- 1101000000100001  lw	r1, r4
  734=>x"1E41",	-- 0001111001000001  mixll	r1, r0, r1
  735=>x"D221",	-- 1101001000100001  sw	r1, r4
  736=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  737=>x"0412",	-- 0000010000010010  inc	r2, r2
  738=>x"061B",	-- 0000011000011011  dec	r3, r3
  739=>x"E398",	-- 1110001110011000  baeq	r3, r6
  740=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop0
  741=>x"D010",	-- 1101000000010000  lw	r0, r2
  742=>x"D021",	-- 1101000000100001  lw	r1, r4
  743=>x"1809",	-- 0001100000001001  mixhh	r1, r1, r0
  744=>x"D221",	-- 1101001000100001  sw	r1, r4
  745=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  746=>x"061B",	-- 0000011000011011  dec	r3, r3
  747=>x"E398",	-- 1110001110011000  baeq	r3, r6
  748=>x"D021",	-- 1101000000100001  lw	r1, r4
  749=>x"1A09",	-- 0001101000001001  mixhl	r1, r1, r0
  750=>x"D221",	-- 1101001000100001  sw	r1, r4
  751=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  752=>x"0412",	-- 0000010000010010  inc	r2, r2
  753=>x"061B",	-- 0000011000011011  dec	r3, r3
  754=>x"E398",	-- 1110001110011000  baeq	r3, r6
  755=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop1
  756=>x"C03D",	-- 1100000000111101  li	r5, 7
  757=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  758=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  759=>x"B5E8",	-- 1011010111101000  brieq	r5, put_sprite_8_aligned
  760=>x"062D",	-- 0000011000101101  dec	r5, r5
  761=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  762=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  763=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  764=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  765=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  766=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  767=>x"8A04",	-- 1000101000000100  brine	r0, put_sprite_8.loop1
  768=>x"D010",	-- 1101000000010000  lw	r0, r2
  769=>x"063F",	-- 0000011000111111  dec	r7, r7
  770=>x"D23A",	-- 1101001000111010  sw	r2, r7
  771=>x"C802",	-- 1100100000000010  li	r2, 0x100
  772=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  773=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  774=>x"D021",	-- 1101000000100001  lw	r1, r4
  775=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  776=>x"2612",	-- 0010011000010010  not	r2, r2
  777=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  778=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  779=>x"D221",	-- 1101001000100001  sw	r1, r4
  780=>x"C0A1",	-- 1100000010100001  li	r1, 20
  781=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  782=>x"D03A",	-- 1101000000111010  lw	r2, r7
  783=>x"043F",	-- 0000010000111111  inc	r7, r7
  784=>x"061B",	-- 0000011000011011  dec	r3, r3
  785=>x"E398",	-- 1110001110011000  baeq	r3, r6
  786=>x"D010",	-- 1101000000010000  lw	r0, r2
  787=>x"063F",	-- 0000011000111111  dec	r7, r7
  788=>x"D23A",	-- 1101001000111010  sw	r2, r7
  789=>x"1E00",	-- 0001111000000000  mixll	r0, r0, r0
  790=>x"C802",	-- 1100100000000010  li	r2, 0x100
  791=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  792=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  793=>x"D021",	-- 1101000000100001  lw	r1, r4
  794=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  795=>x"2612",	-- 0010011000010010  not	r2, r2
  796=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  797=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  798=>x"D221",	-- 1101001000100001  sw	r1, r4
  799=>x"C0A1",	-- 1100000010100001  li	r1, 20
  800=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  801=>x"D03A",	-- 1101000000111010  lw	r2, r7
  802=>x"043F",	-- 0000010000111111  inc	r7, r7
  803=>x"0412",	-- 0000010000010010  inc	r2, r2
  804=>x"061B",	-- 0000011000011011  dec	r3, r3
  805=>x"E398",	-- 1110001110011000  baeq	r3, r6
  806=>x"B683",	-- 1011011010000011  bri	-, put_sprite_8.loop0
  807=>x"D010",	-- 1101000000010000  lw	r0, r2
  808=>x"063F",	-- 0000011000111111  dec	r7, r7
  809=>x"D23A",	-- 1101001000111010  sw	r2, r7
  810=>x"063F",	-- 0000011000111111  dec	r7, r7
  811=>x"D23B",	-- 1101001000111011  sw	r3, r7
  812=>x"C802",	-- 1100100000000010  li	r2, 0x100
  813=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  814=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  815=>x"2080",	-- 0010000010000000  and	r0, r0, r2
  816=>x"D021",	-- 1101000000100001  lw	r1, r4
  817=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
  818=>x"261B",	-- 0010011000011011  not	r3, r3
  819=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  820=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
  821=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  822=>x"D221",	-- 1101001000100001  sw	r1, r4
  823=>x"0424",	-- 0000010000100100  inc	r4, r4
  824=>x"D021",	-- 1101000000100001  lw	r1, r4
  825=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  826=>x"261B",	-- 0010011000011011  not	r3, r3
  827=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  828=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
  829=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  830=>x"D221",	-- 1101001000100001  sw	r1, r4
  831=>x"C099",	-- 1100000010011001  li	r1, 19
  832=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  833=>x"D03B",	-- 1101000000111011  lw	r3, r7
  834=>x"043F",	-- 0000010000111111  inc	r7, r7
  835=>x"D03A",	-- 1101000000111010  lw	r2, r7
  836=>x"043F",	-- 0000010000111111  inc	r7, r7
  837=>x"061B",	-- 0000011000011011  dec	r3, r3
  838=>x"E398",	-- 1110001110011000  baeq	r3, r6
  839=>x"D010",	-- 1101000000010000  lw	r0, r2
  840=>x"4E00",	-- 0100111000000000  shl	r0, r0, 7
  841=>x"063F",	-- 0000011000111111  dec	r7, r7
  842=>x"D23A",	-- 1101001000111010  sw	r2, r7
  843=>x"063F",	-- 0000011000111111  dec	r7, r7
  844=>x"D23B",	-- 1101001000111011  sw	r3, r7
  845=>x"C802",	-- 1100100000000010  li	r2, 0x100
  846=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  847=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  848=>x"2080",	-- 0010000010000000  and	r0, r0, r2
  849=>x"D021",	-- 1101000000100001  lw	r1, r4
  850=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
  851=>x"261B",	-- 0010011000011011  not	r3, r3
  852=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  853=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
  854=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  855=>x"D221",	-- 1101001000100001  sw	r1, r4
  856=>x"0424",	-- 0000010000100100  inc	r4, r4
  857=>x"D021",	-- 1101000000100001  lw	r1, r4
  858=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  859=>x"261B",	-- 0010011000011011  not	r3, r3
  860=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  861=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
  862=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  863=>x"D221",	-- 1101001000100001  sw	r1, r4
  864=>x"C099",	-- 1100000010011001  li	r1, 19
  865=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  866=>x"D03B",	-- 1101000000111011  lw	r3, r7
  867=>x"043F",	-- 0000010000111111  inc	r7, r7
  868=>x"D03A",	-- 1101000000111010  lw	r2, r7
  869=>x"043F",	-- 0000010000111111  inc	r7, r7
  870=>x"0412",	-- 0000010000010010  inc	r2, r2
  871=>x"061B",	-- 0000011000011011  dec	r3, r3
  872=>x"E398",	-- 1110001110011000  baeq	r3, r6
  873=>x"AF83",	-- 1010111110000011  bri	-, put_sprite_8.loop1
    others => x"0000"
    );
begin
  process(CLK)
  begin
    if (CLK'event AND CLK='1') then
      D <= m(to_integer(unsigned(AD)));
    end if;
  end process;
end Behavioral;
