----------------------------------------------------------------------------------
--
-- File retrieved, on 07/02/2010, from :
-- http://sebastien-viardot.imag.fr/Enseignements/Archi1A2s/sources/ROMPROG.vhd
--
-- Slightly altered to get rid of vendor-specific packages and adjust formatting
-- Now auto-filled by asrom script
--
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROMPROG is
  Port ( AD : in  STD_LOGIC_VECTOR (12 downto 0);
         D : out  STD_LOGIC_VECTOR (15 downto 0);
         CLK : in STD_LOGIC);
end ROMPROG;

architecture Behavioral of ROMPROG is
  constant low_address: natural := 0;
  constant high_address: natural := 8192;
  subtype octet is std_logic_vector( 15 downto 0 );
  type zone_memoire is
    array (natural range low_address to high_address-1) of octet;
  constant m: zone_memoire:= (
    0=>x"FFF7",	-- 1111111111110111  liw	r7, IRQ_mask
    1=>x"2000",	-- 0010000000000000  
    2=>x"F8C0",	-- 1111100011000000  bai	-, os_init
    3=>x"0100",	-- 0000000100000000  
   16=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_ack
   17=>x"2002",	-- 0010000000000010  
   18=>x"D001",	-- 1101000000000001  lw	r1, r0
   19=>x"F54A",	-- 1111010101001010  bspl	r2, r1, 5
   20=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_error
   21=>x"0050",	-- 0000000001010000  
   22=>x"F4CA",	-- 1111010011001010  bspl	r2, r1, 3
   23=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_kbd
   24=>x"0060",	-- 0000000001100000  
   25=>x"F40A",	-- 1111010000001010  bspl	r2, r1, 0
   26=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_tmr
   27=>x"0040",	-- 0000000001000000  
   28=>x"D201",	-- 1101001000000001  sw	r1, r0
   29=>x"FFFE",	-- 1111111111111110  reti
   64=>x"263F",	-- 0010011000111111  not r7, r7
   65=>x"D7C0",	-- 1101011111000000  out	r7
   66=>x"E383",	-- 1110001110000011  ba	-, r6
   80=>x"25FF",	-- 0010010111111111  xor	r7, r7, r7
   81=>x"D7C0",	-- 1101011111000000  out	r7
   82=>x"E383",	-- 1110001110000011  ba	-, r6
   96=>x"FFF2",	-- 1111111111110010  liw	r2, PS2_rx
   97=>x"2004",	-- 0010000000000100  
   98=>x"D012",	-- 1101000000010010  lw	r2, r2
   99=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map + 8
  100=>x"16C8",	-- 0001011011001000  
  101=>x"D01B",	-- 1101000000011011  lw	r3, r3
  102=>x"1EBF",	-- 0001111010111111  mixll	r7, r7, r2
  103=>x"C784",	-- 1100011110000100  li	r4, 0xF0
  104=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  105=>x"8C60",	-- 1000110001100000  brieq	r4, int_kbd.release
  106=>x"C704",	-- 1100011100000100  li	r4, 0xE0
  107=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  108=>x"8A20",	-- 1000101000100000  brieq	r4, int_kbd.extended
  109=>x"FFF5",	-- 1111111111110101  liw	r5, rand_seed
  110=>x"16C8",	-- 0001011011001000  
  111=>x"D02C",	-- 1101000000101100  lw	r4, r5
  112=>x"24A4",	-- 0010010010100100  xor	r4, r4, r2
  113=>x"D22C",	-- 1101001000101100  sw	r4, r5
  114=>x"FFF5",	-- 1111111111110101  liw	r5, paper_keys - 1
  115=>x"16CF",	-- 0001011011001111  
  116=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  117=>x"80E0",	-- 1000000011100000  brieq	r4, $+3
  118=>x"FFF5",	-- 1111111111110101  liw	r5, paper_keys + 11 - 1
  119=>x"16DA",	-- 0001011011011010  
  120=>x"042D",	-- 0000010000101101  inc	r5, r5
  121=>x"D02C",	-- 1101000000101100  lw	r4, r5
  122=>x"8560",	-- 1000010101100000  brieq	r4, scan_code_mismatch
  123=>x"6E24",	-- 0110111000100100  shr	r4, r4, 7
  124=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  125=>x"BEE4",	-- 1011111011100100  brine	r4, scan_code_loop
  126=>x"D02A",	-- 1101000000101010  lw	r2, r5
  127=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  128=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  129=>x"741B",	-- 0111010000011011  shr	r3, r3, 10
  130=>x"C00D",	-- 1100000000001101  li	r5, 1
  131=>x"0612",	-- 0000011000010010  dec	r2, r2
  132=>x"3AAA",	-- 0011101010101010  rrl	r2, r5, r2
  133=>x"FFF5",	-- 1111111111110101  liw	r5, key_press_map
  134=>x"16C0",	-- 0001011011000000  
  135=>x"08ED",	-- 0000100011101101  add	r5, r5, r3
  136=>x"D02B",	-- 1101000000101011  lw	r3, r5
  137=>x"80E4",	-- 1000000011100100  brine	r4, scan_code_release
  138=>x"229B",	-- 0010001010011011  or	r3, r3, r2
  139=>x"80C3",	-- 1000000011000011  bri	-, scan_code_notify
  140=>x"2612",	-- 0010011000010010  not	r2, r2
  141=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  142=>x"D22B",	-- 1101001000101011  sw	r3, r5
  143=>x"C003",	-- 1100000000000011  li	r3, 0
  144=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  145=>x"16C8",	-- 0001011011001000  
  146=>x"D223",	-- 1101001000100011  sw	r3, r4
  147=>x"E383",	-- 1110001110000011  ba	-, r6
  148=>x"C014",	-- 1100000000010100  li	r4, 2
  149=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  150=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  151=>x"16C8",	-- 0001011011001000  
  152=>x"D223",	-- 1101001000100011  sw	r3, r4
  153=>x"E383",	-- 1110001110000011  ba	-, r6
  154=>x"C00C",	-- 1100000000001100  li	r4, 1
  155=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  156=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  157=>x"16C8",	-- 0001011011001000  
  158=>x"D223",	-- 1101001000100011  sw	r3, r4
  159=>x"E383",	-- 1110001110000011  ba	-, r6
  256=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_mask
  257=>x"2000",	-- 0010000000000000  
  258=>x"C0C9",	-- 1100000011001001  li	r1, 0x19
  259=>x"D201",	-- 1101001000000001  sw	r1, r0
  260=>x"0400",	-- 0000010000000000  inc	r0, r0
  261=>x"CFF9",	-- 1100111111111001  li	r1, -1
  262=>x"D201",	-- 1101001000000001  sw	r1, r0
  263=>x"C03A",	-- 1100000000111010  li	r2, 7
  264=>x"0880",	-- 0000100010000000  add	r0, r0, r2
  265=>x"C0EA",	-- 1100000011101010  li	r2, 0x1D
  266=>x"D202",	-- 1101001000000010  sw	r2, r0
  267=>x"0400",	-- 0000010000000000  inc	r0, r0
  268=>x"C07A",	-- 1100000001111010  li	r2, 15
  269=>x"D202",	-- 1101001000000010  sw	r2, r0
  270=>x"0400",	-- 0000010000000000  inc	r0, r0
  271=>x"C0DA",	-- 1100000011011010  li	r2, 0x1B
  272=>x"D202",	-- 1101001000000010  sw	r2, r0
  273=>x"0400",	-- 0000010000000000  inc	r0, r0
  274=>x"FFF2",	-- 1111111111110010  liw	r2, 817
  275=>x"0331",	-- 0000001100110001  
  276=>x"D202",	-- 1101001000000010  sw	r2, r0
  277=>x"FFF0",	-- 1111111111110000  liw	r0, key_press_map
  278=>x"16C0",	-- 0001011011000000  
  279=>x"C001",	-- 1100000000000001  li	r1, 0
  280=>x"C042",	-- 1100000001000010  li	r2, 8
  281=>x"D201",	-- 1101001000000001  sw	r1, r0
  282=>x"0400",	-- 0000010000000000  inc	r0, r0
  283=>x"0612",	-- 0000011000010010  dec	r2, r2
  284=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  285=>x"8083",	-- 1000000010000011  bri	-, PaperGameStart
  286=>x"8003",	-- 1000000000000011  bri	-, PaperMenuLoop
  287=>x"FFF0",	-- 1111111111110000  liw	r0, paper_score
  288=>x"16C9",	-- 0001011011001001  
  289=>x"C001",	-- 1100000000000001  li	r1, 0
  290=>x"D201",	-- 1101001000000001  sw	r1, r0
  291=>x"FFF0",	-- 1111111111110000  liw	r0, paper_dir
  292=>x"179C",	-- 0001011110011100  
  293=>x"C001",	-- 1100000000000001  li	r1, 0
  294=>x"D201",	-- 1101001000000001  sw	r1, r0
  295=>x"0400",	-- 0000010000000000  inc	r0, r0
  296=>x"FFF1",	-- 1111111111110001  liw	r1, 152 * 8
  297=>x"04C0",	-- 0000010011000000  
  298=>x"D201",	-- 1101001000000001  sw	r1, r0
  299=>x"0400",	-- 0000010000000000  inc	r0, r0
  300=>x"C001",	-- 1100000000000001  li	r1, 0
  301=>x"D201",	-- 1101001000000001  sw	r1, r0
  302=>x"0400",	-- 0000010000000000  inc	r0, r0
  303=>x"FFF1",	-- 1111111111110001  liw	r1, 128 * 8
  304=>x"0400",	-- 0000010000000000  
  305=>x"D201",	-- 1101001000000001  sw	r1, r0
  306=>x"0400",	-- 0000010000000000  inc	r0, r0
  307=>x"C001",	-- 1100000000000001  li	r1, 0
  308=>x"D201",	-- 1101001000000001  sw	r1, r0
  309=>x"0400",	-- 0000010000000000  inc	r0, r0
  310=>x"C0B9",	-- 1100000010111001  li	r1, 23
  311=>x"D201",	-- 1101001000000001  sw	r1, r0
  312=>x"0400",	-- 0000010000000000  inc	r0, r0
  313=>x"C011",	-- 1100000000010001  li	r1, 2
  314=>x"D201",	-- 1101001000000001  sw	r1, r0
  315=>x"0400",	-- 0000010000000000  inc	r0, r0
  316=>x"FFF0",	-- 1111111111110000  liw	r0, paper_tilemap
  317=>x"17B0",	-- 0001011110110000  
  318=>x"C001",	-- 1100000000000001  li	r1, 0
  319=>x"C0C2",	-- 1100000011000010  li	r2, 6*4
  320=>x"D201",	-- 1101001000000001  sw	r1, r0
  321=>x"0400",	-- 0000010000000000  inc	r0, r0
  322=>x"0612",	-- 0000011000010010  dec	r2, r2
  323=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  324=>x"C000",	-- 1100000000000000  li	r0, 0
  325=>x"CFF9",	-- 1100111111111001  li	r1, -1
  326=>x"C0A2",	-- 1100000010100010  li	r2, 20
  327=>x"D201",	-- 1101001000000001  sw	r1, r0
  328=>x"0400",	-- 0000010000000000  inc	r0, r0
  329=>x"0612",	-- 0000011000010010  dec	r2, r2
  330=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  331=>x"C001",	-- 1100000000000001  li	r1, 0
  332=>x"FFF2",	-- 1111111111110010  liw	r2, 18*20
  333=>x"0168",	-- 0000000101101000  
  334=>x"D201",	-- 1101001000000001  sw	r1, r0
  335=>x"0400",	-- 0000010000000000  inc	r0, r0
  336=>x"0612",	-- 0000011000010010  dec	r2, r2
  337=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  338=>x"CFF9",	-- 1100111111111001  li	r1, -1
  339=>x"C0A2",	-- 1100000010100010  li	r2, 20
  340=>x"D201",	-- 1101001000000001  sw	r1, r0
  341=>x"0400",	-- 0000010000000000  inc	r0, r0
  342=>x"0612",	-- 0000011000010010  dec	r2, r2
  343=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  344=>x"C020",	-- 1100000000100000  li	r0, 4
  345=>x"C029",	-- 1100000000101001  li	r1, 5
  346=>x"FFF2",	-- 1111111111110010  liw	r2, paper_title
  347=>x"17A4",	-- 0001011110100100  
  348=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  349=>x"02AB",	-- 0000001010101011  
  350=>x"C090",	-- 1100000010010000  li	r0, 18
  351=>x"C029",	-- 1100000000101001  li	r1, 5
  352=>x"FFF2",	-- 1111111111110010  liw	r2, paper_score
  353=>x"16C9",	-- 0001011011001001  
  354=>x"D012",	-- 1101000000010010  lw	r2, r2
  355=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum
  356=>x"02DA",	-- 0000001011011010  
  357=>x"C778",	-- 1100011101111000  li	r0, 239
  358=>x"C009",	-- 1100000000001001  li	r1, 1
  359=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud
  360=>x"1780",	-- 0001011110000000  
  361=>x"C043",	-- 1100000001000011  li	r3, 8
  362=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  363=>x"03B3",	-- 0000001110110011  
  364=>x"C0F8",	-- 1100000011111000  li	r0, 31
  365=>x"C009",	-- 1100000000001001  li	r1, 1
  366=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  367=>x"17A0",	-- 0001011110100000  
  368=>x"D012",	-- 1101000000010010  lw	r2, r2
  369=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum
  370=>x"02DA",	-- 0000001011011010  
  371=>x"C120",	-- 1100000100100000  li	r0, 36
  372=>x"C009",	-- 1100000000001001  li	r1, 1
  373=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  374=>x"17AA",	-- 0001011110101010  
  375=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  376=>x"02AB",	-- 0000001010101011  
  377=>x"C778",	-- 1100011101111000  li	r0, 239
  378=>x"C051",	-- 1100000001010001  li	r1, 10
  379=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud + 8
  380=>x"1788",	-- 0001011110001000  
  381=>x"C043",	-- 1100000001000011  li	r3, 8
  382=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  383=>x"03B3",	-- 0000001110110011  
  384=>x"C0F8",	-- 1100000011111000  li	r0, 31
  385=>x"C051",	-- 1100000001010001  li	r1, 10
  386=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed + 1
  387=>x"17A1",	-- 0001011110100001  
  388=>x"D012",	-- 1101000000010010  lw	r2, r2
  389=>x"6412",	-- 0110010000010010  shr	r2, r2, 2
  390=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum
  391=>x"02DA",	-- 0000001011011010  
  392=>x"C120",	-- 1100000100100000  li	r0, 36
  393=>x"C051",	-- 1100000001010001  li	r1, 10
  394=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  395=>x"17AA",	-- 0001011110101010  
  396=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  397=>x"02AB",	-- 0000001010101011  
  398=>x"FFF0",	-- 1111111111110000  liw	r0, 20*20
  399=>x"0190",	-- 0000000110010000  
  400=>x"C001",	-- 1100000000000001  li	r1, 0
  401=>x"FFF2",	-- 1111111111110010  liw	r2, 220*20
  402=>x"1130",	-- 0001000100110000  
  403=>x"D201",	-- 1101001000000001  sw	r1, r0
  404=>x"0400",	-- 0000010000000000  inc	r0, r0
  405=>x"0612",	-- 0000011000010010  dec	r2, r2
  406=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  407=>x"FFF5",	-- 1111111111110101  liw	r5, paper_tilemap
  408=>x"17B0",	-- 0001011110110000  
  409=>x"D02C",	-- 1101000000101100  lw	r4, r5
  410=>x"042D",	-- 0000010000101101  inc	r5, r5
  411=>x"8960",	-- 1000100101100000  brieq	r4, PaperGameTileSkip
  412=>x"063F",	-- 0000011000111111  dec	r7, r7
  413=>x"D23D",	-- 1101001000111101  sw	r5, r7
  414=>x"FFF3",	-- 1111111111110011  liw	r3, paper_tilemap
  415=>x"17B0",	-- 0001011110110000  
  416=>x"0AEB",	-- 0000101011101011  sub	r3, r5, r3
  417=>x"6E20",	-- 0110111000100000  shr	r0, r4, 7
  418=>x"6219",	-- 0110001000011001  shr	r1, r3, 1
  419=>x"4809",	-- 0100100000001001  shl	r1, r1, 4
  420=>x"C19A",	-- 1100000110011010  li	r2, 51
  421=>x"0889",	-- 0000100010001001  add	r1, r1, r2
  422=>x"FFF2",	-- 1111111111110010  liw	r2, paper_pos + 1
  423=>x"179E",	-- 0001011110011110  
  424=>x"D012",	-- 1101000000010010  lw	r2, r2
  425=>x"6412",	-- 0110010000010010  shr	r2, r2, 2
  426=>x"C0FB",	-- 1100000011111011  li	r3, 31
  427=>x"20D2",	-- 0010000011010010  and	r2, r2, r3
  428=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  429=>x"4E24",	-- 0100111000100100  shl	r4, r4, 7
  430=>x"6E24",	-- 0110111000100100  shr	r4, r4, 7
  431=>x"C00B",	-- 1100000000001011  li	r3, 1
  432=>x"FB06",	-- 1111101100000110  bailne	r0, r6, put_tile
  433=>x"027B",	-- 0000001001111011  
  434=>x"81E0",	-- 1000000111100000  brieq	r4, PaperGameSegmentSkip
  436=>x"C013",	-- 1100000000010011  li	r3, 2
  437=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_tile
  438=>x"027B",	-- 0000001001111011  
  439=>x"0624",	-- 0000011000100100  dec	r4, r4
  440=>x"BF64",	-- 1011111101100100  brine	r4, PaperGameSegmentLoop
  441=>x"C003",	-- 1100000000000011  li	r3, 0
  442=>x"C144",	-- 1100000101000100  li	r4, 40
  443=>x"0B04",	-- 0000101100000100  sub	r4, r0, r4
  444=>x"FB66",	-- 1111101101100110  baillt	r4, r6, put_tile
  445=>x"027B",	-- 0000001001111011  
  446=>x"D03D",	-- 1101000000111101  lw	r5, r7
  447=>x"043F",	-- 0000010000111111  inc	r7, r7
  448=>x"FFF4",	-- 1111111111110100  liw r4, paper_tilemap + 24
  449=>x"17C8",	-- 0001011111001000  
  450=>x"0B2C",	-- 0000101100101100  sub	r4, r5, r4
  451=>x"B5A5",	-- 1011010110100101  brilt	r4, PaperGameTileLoop
  452=>x"FFF3",	-- 1111111111110011  liw	r3, paper_speed
  453=>x"17A0",	-- 0001011110100000  
  454=>x"D01B",	-- 1101000000011011  lw	r3, r3
  455=>x"CF04",	-- 1100111100000100  li	r4, 0x1E0
  456=>x"211C",	-- 0010000100011100  and	r4, r3, r4
  457=>x"FFF3",	-- 1111111111110011  liw	r3, paper_pos
  458=>x"179D",	-- 0001011110011101  
  459=>x"D018",	-- 1101000000011000  lw	r0, r3
  460=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  461=>x"FFF2",	-- 1111111111110010  liw	r2, paper_sprites
  462=>x"1720",	-- 0001011100100000  
  463=>x"0912",	-- 0000100100010010  add	r2, r2, r4
  464=>x"C161",	-- 1100000101100001  li	r1, 44
  465=>x"C083",	-- 1100000010000011  li	r3, 16
  466=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_16_masked
  467=>x"034B",	-- 0000001101001011  
  468=>x"902C",	-- 1001000000101100  brine	r5, PaperGameFail
  470=>x"C010",	-- 1100000000010000  li	r0, 2
  471=>x"C001",	-- 1100000000000001  li	r1, 0
  472=>x"8043",	-- 1000000001000011  bri	-, $+1
  473=>x"0609",	-- 0000011000001001  dec	r1, r1
  474=>x"BF8C",	-- 1011111110001100  brine	r1, $-2
  475=>x"0600",	-- 0000011000000000  dec	r0, r0
  476=>x"BEC4",	-- 1011111011000100  brine	r0, $-5
  477=>x"FFF2",	-- 1111111111110010  liw	r2, paper_pos
  478=>x"179D",	-- 0001011110011101  
  479=>x"FFF3",	-- 1111111111110011  liw	r3, paper_speed
  480=>x"17A0",	-- 0001011110100000  
  481=>x"D010",	-- 1101000000010000  lw	r0, r2
  482=>x"D019",	-- 1101000000011001  lw	r1, r3
  483=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  484=>x"8C05",	-- 1000110000000101  brilt	r0, PaperGameFail
  485=>x"FFF4",	-- 1111111111110100  liw	r4, 304*8
  486=>x"0980",	-- 0000100110000000  
  487=>x"0B04",	-- 0000101100000100  sub	r4, r0, r4
  488=>x"8B21",	-- 1000101100100001  brige	r4, PaperGameFail
  489=>x"D210",	-- 1101001000010000  sw	r0, r2
  490=>x"0412",	-- 0000010000010010  inc	r2, r2
  491=>x"041B",	-- 0000010000011011  inc	r3, r3
  492=>x"D010",	-- 1101000000010000  lw	r0, r2
  493=>x"D019",	-- 1101000000011001  lw	r1, r3
  494=>x"C7FC",	-- 1100011111111100  li	r4, 0xFF
  495=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  496=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  497=>x"2101",	-- 0010000100000001  and	r1, r0, r4
  498=>x"D211",	-- 1101001000010001  sw	r1, r2
  499=>x"2624",	-- 0010011000100100  not	r4, r4
  500=>x"2100",	-- 0010000100000000  and	r0, r0, r4
  501=>x"FB06",	-- 1111101100000110  bailne	r0, r6, PaperMapScroll
  502=>x"0236",	-- 0000001000110110  
  503=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  504=>x"16C0",	-- 0001011011000000  
  505=>x"D01B",	-- 1101000000011011  lw	r3, r3
  506=>x"F818",	-- 1111100000011000  baieq	r3, PaperGameRedraw
  507=>x"0144",	-- 0000000101000100  
  508=>x"F55C",	-- 1111010101011100  bspl	r4, r3, 5
  509=>x"8A24",	-- 1000101000100100  brine	r4, PaperGameQuit
  510=>x"F51C",	-- 1111010100011100  bspl	r4, r3, 4
  511=>x"89E4",	-- 1000100111100100  brine	r4, PaperGamePause
  512=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  513=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveUp
  514=>x"F49C",	-- 1111010010011100  bspl	r4, r3, 2
  515=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveDOWN
  516=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  517=>x"81A0",	-- 1000000110100000  brieq	r4, PaperNoMoveLEFT
  518=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  519=>x"17A0",	-- 0001011110100000  
  520=>x"D010",	-- 1101000000010000  lw	r0, r2
  521=>x"0600",	-- 0000011000000000  dec	r0, r0
  522=>x"D210",	-- 1101001000010000  sw	r0, r2
  523=>x"F4DC",	-- 1111010011011100  bspl	r4, r3, 3
  524=>x"81A0",	-- 1000000110100000  brieq	r4, PaperNoMoveRIGHT
  525=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  526=>x"17A0",	-- 0001011110100000  
  527=>x"D010",	-- 1101000000010000  lw	r0, r2
  528=>x"0400",	-- 0000010000000000  inc	r0, r0
  529=>x"D210",	-- 1101001000010000  sw	r0, r2
  530=>x"F8C0",	-- 1111100011000000  bai	-, PaperGameRedraw
  531=>x"0144",	-- 0000000101000100  
  532=>x"C000",	-- 1100000000000000  li	r0, 0
  533=>x"FFF2",	-- 1111111111110010  liw	r2, 240*20
  534=>x"12C0",	-- 0001001011000000  
  535=>x"D001",	-- 1101000000000001  lw	r1, r0
  536=>x"2609",	-- 0010011000001001  not	r1, r1
  537=>x"D201",	-- 1101001000000001  sw	r1, r0
  538=>x"0400",	-- 0000010000000000  inc	r0, r0
  539=>x"0612",	-- 0000011000010010  dec	r2, r2
  540=>x"BED4",	-- 1011111011010100  brine	r2, $-5
  541=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  542=>x"16C0",	-- 0001011011000000  
  543=>x"D01A",	-- 1101000000011010  lw	r2, r3
  544=>x"BFD4",	-- 1011111111010100  brine	r2, $-1
  545=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  546=>x"16C0",	-- 0001011011000000  
  547=>x"D01A",	-- 1101000000011010  lw	r2, r3
  548=>x"BFD0",	-- 1011111111010000  brieq	r2, $-1
  549=>x"FFFF",	-- 1111111111111111  reset
  550=>x"C080",	-- 1100000010000000  li	r0, 16
  551=>x"C0C1",	-- 1100000011000001  li	r1, 24
  552=>x"FFF2",	-- 1111111111110010  liw	r2, paper_pause
  553=>x"17C8",	-- 0001011111001000  
  554=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  555=>x"02AB",	-- 0000001010101011  
  556=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  557=>x"16C0",	-- 0001011011000000  
  558=>x"D01A",	-- 1101000000011010  lw	r2, r3
  559=>x"BFD4",	-- 1011111111010100  brine	r2, $-1
  560=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  561=>x"16C0",	-- 0001011011000000  
  562=>x"D01A",	-- 1101000000011010  lw	r2, r3
  563=>x"BFD0",	-- 1011111111010000  brieq	r2, $-1
  564=>x"F8C0",	-- 1111100011000000  bai	-, PaperGameRedraw
  565=>x"0144",	-- 0000000101000100  
  566=>x"FFF0",	-- 1111111111110000  liw	r0, paper_tilemap
  567=>x"17B0",	-- 0001011110110000  
  568=>x"C021",	-- 1100000000100001  li	r1, 4
  569=>x"0841",	-- 0000100001000001  add	r1, r0, r1
  570=>x"C0A2",	-- 1100000010100010  li	r2, 5*4
  571=>x"D00B",	-- 1101000000001011  lw	r3, r1
  572=>x"D203",	-- 1101001000000011  sw	r3, r0
  573=>x"0400",	-- 0000010000000000  inc	r0, r0
  574=>x"0409",	-- 0000010000001001  inc	r1, r1
  575=>x"0612",	-- 0000011000010010  dec	r2, r2
  576=>x"BED4",	-- 1011111011010100  brine	r2, PaperGameScrollLoop
  577=>x"063F",	-- 0000011000111111  dec	r7, r7
  578=>x"D23E",	-- 1101001000111110  sw	r6, r7
  579=>x"FAC6",	-- 1111101011000110  bail	-, r6, rand16
  580=>x"0269",	-- 0000001001101001  
  581=>x"FFF2",	-- 1111111111110010  liw	r2, 0x7777
  582=>x"7777",	-- 0111011101110111  
  583=>x"208A",	-- 0010000010001010  and	r2, r1, r2
  584=>x"6613",	-- 0110011000010011  shr	r3, r2, 3
  585=>x"C87C",	-- 1100100001111100  li	r4, 0x10F
  586=>x"211B",	-- 0010000100011011  and	r3, r3, r4
  587=>x"D201",	-- 1101001000000001  sw	r1, r0
  588=>x"0400",	-- 0000010000000000  inc	r0, r0
  589=>x"6E14",	-- 0110111000010100  shr	r4, r2, 7
  590=>x"C07D",	-- 1100000001111101  li	r5, 0x0F
  591=>x"2164",	-- 0010000101100100  and	r4, r4, r5
  592=>x"0424",	-- 0000010000100100  inc	r4, r4
  593=>x"0424",	-- 0000010000100100  inc	r4, r4
  594=>x"0424",	-- 0000010000100100  inc	r4, r4
  595=>x"4E24",	-- 0100111000100100  shl	r4, r4, 7
  596=>x"08E3",	-- 0000100011100011  add	r3, r4, r3
  597=>x"2152",	-- 0010000101010010  and	r2, r2, r5
  598=>x"095B",	-- 0000100101011011  add	r3, r3, r5
  599=>x"D201",	-- 1101001000000001  sw	r1, r0
  600=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed + 1
  601=>x"17A1",	-- 0001011110100001  
  602=>x"D011",	-- 1101000000010001  lw	r1, r2
  603=>x"0409",	-- 0000010000001001  inc	r1, r1
  604=>x"D211",	-- 1101001000010001  sw	r1, r2
  605=>x"FFF2",	-- 1111111111110010  liw	r2, paper_score
  606=>x"16C9",	-- 0001011011001001  
  607=>x"D011",	-- 1101000000010001  lw	r1, r2
  608=>x"0409",	-- 0000010000001001  inc	r1, r1
  609=>x"D211",	-- 1101001000010001  sw	r1, r2
  610=>x"D03E",	-- 1101000000111110  lw	r6, r7
  611=>x"043F",	-- 0000010000111111  inc	r7, r7
  612=>x"E383",	-- 1110001110000011  ba	-, r6
  613=>x"FFF2",	-- 1111111111110010  liw	r2, rand_seed
  614=>x"16C8",	-- 0001011011001000  
  615=>x"D210",	-- 1101001000010000  sw	r0, r2
  616=>x"E383",	-- 1110001110000011  ba	-, r6
  617=>x"FFF2",	-- 1111111111110010  liw	r2, rand_seed
  618=>x"16C8",	-- 0001011011001000  
  619=>x"D013",	-- 1101000000010011  lw	r3, r2
  620=>x"C7EC",	-- 1100011111101100  li	r4, 253
  621=>x"1F19",	-- 0001111100011001  mixll	r1, r3, r4
  622=>x"18E4",	-- 0001100011100100  mixhh	r4, r4, r3
  623=>x"C002",	-- 1100000000000010  li	r2, 0
  624=>x"0AC9",	-- 0000101011001001  sub	r1, r1, r3
  625=>x"0EA4",	-- 0000111010100100  sbc	r4, r4, r2
  626=>x"0EC9",	-- 0000111011001001  sbc	r1, r1, r3
  627=>x"0EA4",	-- 0000111010100100  sbc	r4, r4, r2
  628=>x"1B13",	-- 0001101100010011  mixhl	r3, r2, r4
  629=>x"0EC9",	-- 0000111011001001  sbc	r1, r1, r3
  630=>x"0C89",	-- 0000110010001001  adc	r1, r1, r2
  631=>x"FFF2",	-- 1111111111110010  liw	r2, rand_seed
  632=>x"16C8",	-- 0001011011001000  
  633=>x"D211",	-- 1101001000010001  sw	r1, r2
  634=>x"E383",	-- 1110001110000011  ba	-, r6
  635=>x"063F",	-- 0000011000111111  dec	r7, r7
  636=>x"D238",	-- 1101001000111000  sw	r0, r7
  637=>x"063F",	-- 0000011000111111  dec	r7, r7
  638=>x"D239",	-- 1101001000111001  sw	r1, r7
  639=>x"063F",	-- 0000011000111111  dec	r7, r7
  640=>x"D23A",	-- 1101001000111010  sw	r2, r7
  641=>x"063F",	-- 0000011000111111  dec	r7, r7
  642=>x"D23B",	-- 1101001000111011  sw	r3, r7
  643=>x"063F",	-- 0000011000111111  dec	r7, r7
  644=>x"D23C",	-- 1101001000111100  sw	r4, r7
  645=>x"063F",	-- 0000011000111111  dec	r7, r7
  646=>x"D23D",	-- 1101001000111101  sw	r5, r7
  647=>x"063F",	-- 0000011000111111  dec	r7, r7
  648=>x"D23E",	-- 1101001000111110  sw	r6, r7
  649=>x"FFF2",	-- 1111111111110010  liw	r2, paper_tiles
  650=>x"1790",	-- 0001011110010000  
  651=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  652=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  653=>x"C043",	-- 1100000001000011  li	r3, 8
  654=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  655=>x"038D",	-- 0000001110001101  
  656=>x"D03E",	-- 1101000000111110  lw	r6, r7
  657=>x"043F",	-- 0000010000111111  inc	r7, r7
  658=>x"D03D",	-- 1101000000111101  lw	r5, r7
  659=>x"043F",	-- 0000010000111111  inc	r7, r7
  660=>x"D03C",	-- 1101000000111100  lw	r4, r7
  661=>x"043F",	-- 0000010000111111  inc	r7, r7
  662=>x"D03B",	-- 1101000000111011  lw	r3, r7
  663=>x"043F",	-- 0000010000111111  inc	r7, r7
  664=>x"D03A",	-- 1101000000111010  lw	r2, r7
  665=>x"043F",	-- 0000010000111111  inc	r7, r7
  666=>x"D039",	-- 1101000000111001  lw	r1, r7
  667=>x"043F",	-- 0000010000111111  inc	r7, r7
  668=>x"D038",	-- 1101000000111000  lw	r0, r7
  669=>x"043F",	-- 0000010000111111  inc	r7, r7
  670=>x"0400",	-- 0000010000000000  inc	r0, r0
  671=>x"E383",	-- 1110001110000011  ba	-, r6
  672=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  673=>x"C084",	-- 1100000010000100  li	r4, 16
  674=>x"0800",	-- 0000100000000000  add	r0, r0, r0
  675=>x"0C49",	-- 0000110001001001  adc	r1, r1, r1
  676=>x"0A8B",	-- 0000101010001011  sub	r3, r1, r2
  677=>x"80DD",	-- 1000000011011101  brilt	r3, div_16_16.skip
  678=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  679=>x"0400",	-- 0000010000000000  inc	r0, r0
  680=>x"0624",	-- 0000011000100100  dec	r4, r4
  681=>x"BE64",	-- 1011111001100100  brine	r4, div_16_16.loop
  682=>x"E383",	-- 1110001110000011  ba	-, r6
  683=>x"063F",	-- 0000011000111111  dec	r7, r7
  684=>x"D23E",	-- 1101001000111110  sw	r6, r7
  685=>x"D013",	-- 1101000000010011  lw	r3, r2
  686=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  687=>x"84D8",	-- 1000010011011000  brieq	r3, puts.end
  688=>x"063F",	-- 0000011000111111  dec	r7, r7
  689=>x"D23A",	-- 1101001000111010  sw	r2, r7
  690=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  691=>x"02C5",	-- 0000001011000101  
  692=>x"D03A",	-- 1101000000111010  lw	r2, r7
  693=>x"043F",	-- 0000010000111111  inc	r7, r7
  694=>x"D013",	-- 1101000000010011  lw	r3, r2
  695=>x"4E1B",	-- 0100111000011011  shl	r3, r3, 7
  696=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  697=>x"8258",	-- 1000001001011000  brieq	r3, puts.end
  698=>x"063F",	-- 0000011000111111  dec	r7, r7
  699=>x"D23A",	-- 1101001000111010  sw	r2, r7
  700=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  701=>x"02C5",	-- 0000001011000101  
  702=>x"D03A",	-- 1101000000111010  lw	r2, r7
  703=>x"043F",	-- 0000010000111111  inc	r7, r7
  704=>x"0412",	-- 0000010000010010  inc	r2, r2
  705=>x"BB03",	-- 1011101100000011  bri	-, puts.loop
  706=>x"D03E",	-- 1101000000111110  lw	r6, r7
  707=>x"043F",	-- 0000010000111111  inc	r7, r7
  708=>x"E383",	-- 1110001110000011  ba	-, r6
  709=>x"063F",	-- 0000011000111111  dec	r7, r7
  710=>x"D23E",	-- 1101001000111110  sw	r6, r7
  711=>x"063F",	-- 0000011000111111  dec	r7, r7
  712=>x"D238",	-- 1101001000111000  sw	r0, r7
  713=>x"063F",	-- 0000011000111111  dec	r7, r7
  714=>x"D239",	-- 1101001000111001  sw	r1, r7
  715=>x"FFF2",	-- 1111111111110010  liw	r2, font_map
  716=>x"12C0",	-- 0001001011000000  
  717=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  718=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  719=>x"C043",	-- 1100000001000011  li	r3, 8
  720=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  721=>x"038D",	-- 0000001110001101  
  722=>x"D039",	-- 1101000000111001  lw	r1, r7
  723=>x"043F",	-- 0000010000111111  inc	r7, r7
  724=>x"D038",	-- 1101000000111000  lw	r0, r7
  725=>x"043F",	-- 0000010000111111  inc	r7, r7
  726=>x"0400",	-- 0000010000000000  inc	r0, r0
  727=>x"D03E",	-- 1101000000111110  lw	r6, r7
  728=>x"043F",	-- 0000010000111111  inc	r7, r7
  729=>x"E383",	-- 1110001110000011  ba	-, r6
  730=>x"063F",	-- 0000011000111111  dec	r7, r7
  731=>x"D23E",	-- 1101001000111110  sw	r6, r7
  732=>x"FFF4",	-- 1111111111110100  liw	r4, 10000
  733=>x"2710",	-- 0010011100010000  
  734=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  735=>x"02ED",	-- 0000001011101101  
  736=>x"FFF4",	-- 1111111111110100  liw	r4, 1000
  737=>x"03E8",	-- 0000001111101000  
  738=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  739=>x"02ED",	-- 0000001011101101  
  740=>x"C324",	-- 1100001100100100  li	r4, 100
  741=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  742=>x"02ED",	-- 0000001011101101  
  743=>x"C054",	-- 1100000001010100  li	r4, 10
  744=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  745=>x"02ED",	-- 0000001011101101  
  746=>x"D03E",	-- 1101000000111110  lw	r6, r7
  747=>x"043F",	-- 0000010000111111  inc	r7, r7
  748=>x"C00C",	-- 1100000000001100  li	r4, 1
  749=>x"C17B",	-- 1100000101111011  li	r3, 0x2F
  750=>x"041B",	-- 0000010000011011  inc	r3, r3
  751=>x"0B12",	-- 0000101100010010  sub	r2, r2, r4
  752=>x"BF91",	-- 1011111110010001  brige	r2, printnum.loop
  753=>x"0912",	-- 0000100100010010  add	r2, r2, r4
  754=>x"063F",	-- 0000011000111111  dec	r7, r7
  755=>x"D23E",	-- 1101001000111110  sw	r6, r7
  756=>x"063F",	-- 0000011000111111  dec	r7, r7
  757=>x"D23A",	-- 1101001000111010  sw	r2, r7
  758=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  759=>x"02C5",	-- 0000001011000101  
  760=>x"D03A",	-- 1101000000111010  lw	r2, r7
  761=>x"043F",	-- 0000010000111111  inc	r7, r7
  762=>x"D03E",	-- 1101000000111110  lw	r6, r7
  763=>x"043F",	-- 0000010000111111  inc	r7, r7
  764=>x"E383",	-- 1110001110000011  ba	-, r6
  765=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  766=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  767=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  768=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  769=>x"C0A0",	-- 1100000010100000  li	r0, 20
  770=>x"0412",	-- 0000010000010010  inc	r2, r2
  771=>x"D011",	-- 1101000000010001  lw	r1, r2
  772=>x"E421",	-- 1110010000100001  exw	r1, r4
  773=>x"0412",	-- 0000010000010010  inc	r2, r2
  774=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  775=>x"061B",	-- 0000011000011011  dec	r3, r3
  776=>x"BE9C",	-- 1011111010011100  brine	r3, put_sprite_16_aligned.loop
  777=>x"C005",	-- 1100000000000101  li	r5, 0
  778=>x"E383",	-- 1110001110000011  ba	-, r6
  779=>x"C07D",	-- 1100000001111101  li	r5, 15
  780=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  781=>x"6600",	-- 0110011000000000  shr	r0, r0, 3
  782=>x"BBE8",	-- 1011101111101000  brieq	r5, put_sprite_16_aligned
  783=>x"062D",	-- 0000011000101101  dec	r5, r5
  784=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  785=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  786=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  787=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  788=>x"063F",	-- 0000011000111111  dec	r7, r7
  789=>x"D23B",	-- 1101001000111011  sw	r3, r7
  790=>x"0412",	-- 0000010000010010  inc	r2, r2
  791=>x"D011",	-- 1101000000010001  lw	r1, r2
  792=>x"CFF8",	-- 1100111111111000  li	r0, -1
  793=>x"3D40",	-- 0011110101000000  rsr	r0, r0, r5
  794=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  795=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  796=>x"D023",	-- 1101000000100011  lw	r3, r4
  797=>x"2600",	-- 0010011000000000  not	r0, r0
  798=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  799=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  800=>x"E421",	-- 1110010000100001  exw	r1, r4
  801=>x"0424",	-- 0000010000100100  inc	r4, r4
  802=>x"D011",	-- 1101000000010001  lw	r1, r2
  803=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  804=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  805=>x"D023",	-- 1101000000100011  lw	r3, r4
  806=>x"2600",	-- 0010011000000000  not	r0, r0
  807=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  808=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  809=>x"E421",	-- 1110010000100001  exw	r1, r4
  810=>x"0412",	-- 0000010000010010  inc	r2, r2
  811=>x"C098",	-- 1100000010011000  li	r0, 19
  812=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  813=>x"D03B",	-- 1101000000111011  lw	r3, r7
  814=>x"043F",	-- 0000010000111111  inc	r7, r7
  815=>x"061B",	-- 0000011000011011  dec	r3, r3
  816=>x"B91C",	-- 1011100100011100  brine	r3, put_sprite_16.loop
  817=>x"C005",	-- 1100000000000101  li	r5, 0
  818=>x"E383",	-- 1110001110000011  ba	-, r6
  819=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  820=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  821=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  822=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  823=>x"C005",	-- 1100000000000101  li	r5, 0
  824=>x"D020",	-- 1101000000100000  lw	r0, r4
  825=>x"D011",	-- 1101000000010001  lw	r1, r2
  826=>x"0412",	-- 0000010000010010  inc	r2, r2
  827=>x"2040",	-- 0010000001000000  and	r0, r0, r1
  828=>x"D011",	-- 1101000000010001  lw	r1, r2
  829=>x"2240",	-- 0010001001000000  or	r0, r0, r1
  830=>x"E420",	-- 1110010000100000  exw	r0, r4
  831=>x"0612",	-- 0000011000010010  dec	r2, r2
  832=>x"D011",	-- 1101000000010001  lw	r1, r2
  833=>x"2609",	-- 0010011000001001  not	r1, r1
  834=>x"0412",	-- 0000010000010010  inc	r2, r2
  835=>x"2040",	-- 0010000001000000  and	r0, r0, r1
  836=>x"222D",	-- 0010001000101101  or	r5, r5, r0
  837=>x"0412",	-- 0000010000010010  inc	r2, r2
  838=>x"C0A0",	-- 1100000010100000  li	r0, 20
  839=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  840=>x"061B",	-- 0000011000011011  dec	r3, r3
  841=>x"AE5C",	-- 1010111001011100  brine	r3, put_sprite_16_aligned.loop
  842=>x"E383",	-- 1110001110000011  ba	-, r6
  843=>x"C07D",	-- 1100000001111101  li	r5, 15
  844=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  845=>x"6600",	-- 0110011000000000  shr	r0, r0, 3
  846=>x"B968",	-- 1011100101101000  brieq	r5, put_sprite_16_masked_aligned
  847=>x"062D",	-- 0000011000101101  dec	r5, r5
  848=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  849=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  850=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  851=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  852=>x"063F",	-- 0000011000111111  dec	r7, r7
  853=>x"D23E",	-- 1101001000111110  sw	r6, r7
  854=>x"102E",	-- 0001000000101110  mova	r6, r5
  855=>x"C005",	-- 1100000000000101  li	r5, 0
  856=>x"063F",	-- 0000011000111111  dec	r7, r7
  857=>x"D23B",	-- 1101001000111011  sw	r3, r7
  858=>x"063F",	-- 0000011000111111  dec	r7, r7
  859=>x"D23D",	-- 1101001000111101  sw	r5, r7
  860=>x"D010",	-- 1101000000010000  lw	r0, r2
  861=>x"3980",	-- 0011100110000000  rrr	r0, r0, r6
  862=>x"0412",	-- 0000010000010010  inc	r2, r2
  863=>x"D011",	-- 1101000000010001  lw	r1, r2
  864=>x"3989",	-- 0011100110001001  rrr	r1, r1, r6
  865=>x"CFFD",	-- 1100111111111101  li	r5, -1
  866=>x"3DAD",	-- 0011110110101101  rsr	r5, r5, r6
  867=>x"2149",	-- 0010000101001001  and	r1, r1, r5
  868=>x"D023",	-- 1101000000100011  lw	r3, r4
  869=>x"262D",	-- 0010011000101101  not	r5, r5
  870=>x"222D",	-- 0010001000101101  or	r5, r5, r0
  871=>x"215B",	-- 0010000101011011  and	r3, r3, r5
  872=>x"225B",	-- 0010001001011011  or	r3, r3, r1
  873=>x"E423",	-- 1110010000100011  exw	r3, r4
  874=>x"262D",	-- 0010011000101101  not	r5, r5
  875=>x"215B",	-- 0010000101011011  and	r3, r3, r5
  876=>x"D03D",	-- 1101000000111101  lw	r5, r7
  877=>x"043F",	-- 0000010000111111  inc	r7, r7
  878=>x"22ED",	-- 0010001011101101  or	r5, r5, r3
  879=>x"0424",	-- 0000010000100100  inc	r4, r4
  880=>x"063F",	-- 0000011000111111  dec	r7, r7
  881=>x"D23D",	-- 1101001000111101  sw	r5, r7
  882=>x"D011",	-- 1101000000010001  lw	r1, r2
  883=>x"3989",	-- 0011100110001001  rrr	r1, r1, r6
  884=>x"CFFD",	-- 1100111111111101  li	r5, -1
  885=>x"3DAD",	-- 0011110110101101  rsr	r5, r5, r6
  886=>x"262D",	-- 0010011000101101  not	r5, r5
  887=>x"2149",	-- 0010000101001001  and	r1, r1, r5
  888=>x"D023",	-- 1101000000100011  lw	r3, r4
  889=>x"262D",	-- 0010011000101101  not	r5, r5
  890=>x"222D",	-- 0010001000101101  or	r5, r5, r0
  891=>x"215B",	-- 0010000101011011  and	r3, r3, r5
  892=>x"225B",	-- 0010001001011011  or	r3, r3, r1
  893=>x"E423",	-- 1110010000100011  exw	r3, r4
  894=>x"262D",	-- 0010011000101101  not	r5, r5
  895=>x"215B",	-- 0010000101011011  and	r3, r3, r5
  896=>x"D03D",	-- 1101000000111101  lw	r5, r7
  897=>x"043F",	-- 0000010000111111  inc	r7, r7
  898=>x"22ED",	-- 0010001011101101  or	r5, r5, r3
  899=>x"0412",	-- 0000010000010010  inc	r2, r2
  900=>x"C098",	-- 1100000010011000  li	r0, 19
  901=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  902=>x"D03B",	-- 1101000000111011  lw	r3, r7
  903=>x"043F",	-- 0000010000111111  inc	r7, r7
  904=>x"061B",	-- 0000011000011011  dec	r3, r3
  905=>x"B3DC",	-- 1011001111011100  brine	r3, put_sprite_16_masked.loop
  906=>x"D03E",	-- 1101000000111110  lw	r6, r7
  907=>x"043F",	-- 0000010000111111  inc	r7, r7
  908=>x"E383",	-- 1110001110000011  ba	-, r6
  909=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  910=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  911=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  912=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  913=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  914=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  915=>x"C0A5",	-- 1100000010100101  li	r5, 20
  916=>x"8404",	-- 1000010000000100  brine	r0, put_sprite_8_aligned.loop1
  917=>x"D010",	-- 1101000000010000  lw	r0, r2
  918=>x"D021",	-- 1101000000100001  lw	r1, r4
  919=>x"1A41",	-- 0001101001000001  mixhl	r1, r0, r1
  920=>x"D221",	-- 1101001000100001  sw	r1, r4
  921=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  922=>x"061B",	-- 0000011000011011  dec	r3, r3
  923=>x"E398",	-- 1110001110011000  baeq	r3, r6
  924=>x"D021",	-- 1101000000100001  lw	r1, r4
  925=>x"1E41",	-- 0001111001000001  mixll	r1, r0, r1
  926=>x"D221",	-- 1101001000100001  sw	r1, r4
  927=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  928=>x"0412",	-- 0000010000010010  inc	r2, r2
  929=>x"061B",	-- 0000011000011011  dec	r3, r3
  930=>x"E398",	-- 1110001110011000  baeq	r3, r6
  931=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop0
  932=>x"D010",	-- 1101000000010000  lw	r0, r2
  933=>x"D021",	-- 1101000000100001  lw	r1, r4
  934=>x"1809",	-- 0001100000001001  mixhh	r1, r1, r0
  935=>x"D221",	-- 1101001000100001  sw	r1, r4
  936=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  937=>x"061B",	-- 0000011000011011  dec	r3, r3
  938=>x"E398",	-- 1110001110011000  baeq	r3, r6
  939=>x"D021",	-- 1101000000100001  lw	r1, r4
  940=>x"1A09",	-- 0001101000001001  mixhl	r1, r1, r0
  941=>x"D221",	-- 1101001000100001  sw	r1, r4
  942=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  943=>x"0412",	-- 0000010000010010  inc	r2, r2
  944=>x"061B",	-- 0000011000011011  dec	r3, r3
  945=>x"E398",	-- 1110001110011000  baeq	r3, r6
  946=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop1
  947=>x"C03D",	-- 1100000000111101  li	r5, 7
  948=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  949=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  950=>x"B5E8",	-- 1011010111101000  brieq	r5, put_sprite_8_aligned
  951=>x"062D",	-- 0000011000101101  dec	r5, r5
  952=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  953=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  954=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  955=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  956=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  957=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  958=>x"8A04",	-- 1000101000000100  brine	r0, put_sprite_8.loop1
  959=>x"D010",	-- 1101000000010000  lw	r0, r2
  960=>x"063F",	-- 0000011000111111  dec	r7, r7
  961=>x"D23A",	-- 1101001000111010  sw	r2, r7
  962=>x"C802",	-- 1100100000000010  li	r2, 0x100
  963=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  964=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  965=>x"D021",	-- 1101000000100001  lw	r1, r4
  966=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  967=>x"2612",	-- 0010011000010010  not	r2, r2
  968=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  969=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  970=>x"D221",	-- 1101001000100001  sw	r1, r4
  971=>x"C0A1",	-- 1100000010100001  li	r1, 20
  972=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  973=>x"D03A",	-- 1101000000111010  lw	r2, r7
  974=>x"043F",	-- 0000010000111111  inc	r7, r7
  975=>x"061B",	-- 0000011000011011  dec	r3, r3
  976=>x"E398",	-- 1110001110011000  baeq	r3, r6
  977=>x"D010",	-- 1101000000010000  lw	r0, r2
  978=>x"063F",	-- 0000011000111111  dec	r7, r7
  979=>x"D23A",	-- 1101001000111010  sw	r2, r7
  980=>x"1E00",	-- 0001111000000000  mixll	r0, r0, r0
  981=>x"C802",	-- 1100100000000010  li	r2, 0x100
  982=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  983=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  984=>x"D021",	-- 1101000000100001  lw	r1, r4
  985=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  986=>x"2612",	-- 0010011000010010  not	r2, r2
  987=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  988=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  989=>x"D221",	-- 1101001000100001  sw	r1, r4
  990=>x"C0A1",	-- 1100000010100001  li	r1, 20
  991=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  992=>x"D03A",	-- 1101000000111010  lw	r2, r7
  993=>x"043F",	-- 0000010000111111  inc	r7, r7
  994=>x"0412",	-- 0000010000010010  inc	r2, r2
  995=>x"061B",	-- 0000011000011011  dec	r3, r3
  996=>x"E398",	-- 1110001110011000  baeq	r3, r6
  997=>x"B683",	-- 1011011010000011  bri	-, put_sprite_8.loop0
  998=>x"D010",	-- 1101000000010000  lw	r0, r2
  999=>x"063F",	-- 0000011000111111  dec	r7, r7
 1000=>x"D23A",	-- 1101001000111010  sw	r2, r7
 1001=>x"063F",	-- 0000011000111111  dec	r7, r7
 1002=>x"D23B",	-- 1101001000111011  sw	r3, r7
 1003=>x"C802",	-- 1100100000000010  li	r2, 0x100
 1004=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
 1005=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
 1006=>x"2080",	-- 0010000010000000  and	r0, r0, r2
 1007=>x"D021",	-- 1101000000100001  lw	r1, r4
 1008=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
 1009=>x"261B",	-- 0010011000011011  not	r3, r3
 1010=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
 1011=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
 1012=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
 1013=>x"D221",	-- 1101001000100001  sw	r1, r4
 1014=>x"0424",	-- 0000010000100100  inc	r4, r4
 1015=>x"D021",	-- 1101000000100001  lw	r1, r4
 1016=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
 1017=>x"261B",	-- 0010011000011011  not	r3, r3
 1018=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
 1019=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
 1020=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
 1021=>x"D221",	-- 1101001000100001  sw	r1, r4
 1022=>x"C099",	-- 1100000010011001  li	r1, 19
 1023=>x"0864",	-- 0000100001100100  add	r4, r4, r1
 1024=>x"D03B",	-- 1101000000111011  lw	r3, r7
 1025=>x"043F",	-- 0000010000111111  inc	r7, r7
 1026=>x"D03A",	-- 1101000000111010  lw	r2, r7
 1027=>x"043F",	-- 0000010000111111  inc	r7, r7
 1028=>x"061B",	-- 0000011000011011  dec	r3, r3
 1029=>x"E398",	-- 1110001110011000  baeq	r3, r6
 1030=>x"D010",	-- 1101000000010000  lw	r0, r2
 1031=>x"4E00",	-- 0100111000000000  shl	r0, r0, 7
 1032=>x"063F",	-- 0000011000111111  dec	r7, r7
 1033=>x"D23A",	-- 1101001000111010  sw	r2, r7
 1034=>x"063F",	-- 0000011000111111  dec	r7, r7
 1035=>x"D23B",	-- 1101001000111011  sw	r3, r7
 1036=>x"C802",	-- 1100100000000010  li	r2, 0x100
 1037=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
 1038=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
 1039=>x"2080",	-- 0010000010000000  and	r0, r0, r2
 1040=>x"D021",	-- 1101000000100001  lw	r1, r4
 1041=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
 1042=>x"261B",	-- 0010011000011011  not	r3, r3
 1043=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
 1044=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
 1045=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
 1046=>x"D221",	-- 1101001000100001  sw	r1, r4
 1047=>x"0424",	-- 0000010000100100  inc	r4, r4
 1048=>x"D021",	-- 1101000000100001  lw	r1, r4
 1049=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
 1050=>x"261B",	-- 0010011000011011  not	r3, r3
 1051=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
 1052=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
 1053=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
 1054=>x"D221",	-- 1101001000100001  sw	r1, r4
 1055=>x"C099",	-- 1100000010011001  li	r1, 19
 1056=>x"0864",	-- 0000100001100100  add	r4, r4, r1
 1057=>x"D03B",	-- 1101000000111011  lw	r3, r7
 1058=>x"043F",	-- 0000010000111111  inc	r7, r7
 1059=>x"D03A",	-- 1101000000111010  lw	r2, r7
 1060=>x"043F",	-- 0000010000111111  inc	r7, r7
 1061=>x"0412",	-- 0000010000010010  inc	r2, r2
 1062=>x"061B",	-- 0000011000011011  dec	r3, r3
 1063=>x"E398",	-- 1110001110011000  baeq	r3, r6
 1064=>x"AF83",	-- 1010111110000011  bri	-, put_sprite_8.loop1
    others => x"0000"
    );
begin
  process(CLK)
  begin
    if (CLK'event AND CLK='1') then
      D <= m(to_integer(unsigned(AD)));
    end if;
  end process;
end Behavioral;
