----------------------------------------------------------------------------------
--
-- File retrieved, on 07/02/2010, from :
-- http://sebastien-viardot.imag.fr/Enseignements/Archi1A2s/sources/ROMPROG.vhd
--
-- Slightly altered to get rid of vendor-specific packages and adjust formatting
-- Now auto-filled by asrom script
--
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROMPROG is
  Port ( AD : in  STD_LOGIC_VECTOR (12 downto 0);
         D : out  STD_LOGIC_VECTOR (15 downto 0);
         CLK : in STD_LOGIC);
end ROMPROG;

architecture Behavioral of ROMPROG is
  constant low_address: natural := 0;
  constant high_address: natural := 8192;
  subtype octet is std_logic_vector( 15 downto 0 );
  type zone_memoire is
    array (natural range low_address to high_address-1) of octet;
  constant m: zone_memoire:= (
    0=>x"FFF7",	-- 1111111111110111  liw	r7, IRQ_mask
    1=>x"2000",	-- 0010000000000000  
    2=>x"F8C0",	-- 1111100011000000  bai	-, os_init
    3=>x"0100",	-- 0000000100000000  
   16=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_ack
   17=>x"2002",	-- 0010000000000010  
   18=>x"D001",	-- 1101000000000001  lw	r1, r0
   19=>x"F54A",	-- 1111010101001010  bspl	r2, r1, 5
   20=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_error
   21=>x"00A0",	-- 0000000010100000  
   22=>x"F4CA",	-- 1111010011001010  bspl	r2, r1, 3
   23=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_kbd
   24=>x"0090",	-- 0000000010010000  
   25=>x"F40A",	-- 1111010000001010  bspl	r2, r1, 0
   26=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_tmr
   27=>x"0080",	-- 0000000010000000  
   28=>x"CFF9",	-- 1100111111111001  li	r1, -1
   29=>x"D201",	-- 1101001000000001  sw	r1, r0
   30=>x"FFFE",	-- 1111111111111110  reti
  128=>x"2624",	-- 0010011000100100  not r4, r4
  129=>x"D700",	-- 1101011100000000  out	r4
  130=>x"E383",	-- 1110001110000011  ba	-, r6
  144=>x"E383",	-- 1110001110000011  ba	-, r6
  160=>x"2524",	-- 0010010100100100  xor	r4, r4, r4
  161=>x"D700",	-- 1101011100000000  out	r4
  162=>x"E383",	-- 1110001110000011  ba	-, r6
  256=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_mask
  257=>x"2000",	-- 0010000000000000  
  258=>x"C0C9",	-- 1100000011001001  li	r1, 0x19
  259=>x"D201",	-- 1101001000000001  sw	r1, r0
  260=>x"0400",	-- 0000010000000000  inc	r0, r0
  261=>x"CFF9",	-- 1100111111111001  li	r1, -1
  262=>x"D201",	-- 1101001000000001  sw	r1, r0
  263=>x"C03A",	-- 1100000000111010  li	r2, 7
  264=>x"0880",	-- 0000100010000000  add	r0, r0, r2
  265=>x"C0EA",	-- 1100000011101010  li	r2, 0x1D
  266=>x"D202",	-- 1101001000000010  sw	r2, r0
  267=>x"0400",	-- 0000010000000000  inc	r0, r0
  268=>x"C07A",	-- 1100000001111010  li	r2, 15
  269=>x"D202",	-- 1101001000000010  sw	r2, r0
  270=>x"FFF0",	-- 1111111111110000  liw	r0, 0x8421
  271=>x"8421",	-- 1000010000100001  
  272=>x"FFF1",	-- 1111111111110001  liw	r1, 0x1234
  273=>x"1234",	-- 0001001000110100  
  274=>x"D640",	-- 1101011001000000  out	r1
  275=>x"E408",	-- 1110010000001000  exw	r0, r1
  276=>x"E408",	-- 1110010000001000  exw	r0, r1
  277=>x"1842",	-- 0001100001000010  mixhh	r2, r0, r1
  278=>x"1A43",	-- 0001101001000011  mixhl	r3, r0, r1
  279=>x"1C44",	-- 0001110001000100  mixlh	r4, r0, r1
  280=>x"1E45",	-- 0001111001000101  mixll	r5, r0, r1
  281=>x"C01E",	-- 1100000000011110  li	r6, 3
  282=>x"3985",	-- 0011100110000101  rrr	r5, r0, r6
  283=>x"3B8D",	-- 0011101110001101  rrl	r5, r1, r6
  284=>x"3D95",	-- 0011110110010101  rsr	r5, r2, r6
  285=>x"3F9D",	-- 0011111110011101  rsl	r5, r3, r6
  286=>x"FC0E",	-- 1111110000001110  mul	r6, r1, r0
  287=>x"C138",	-- 1100000100111000  li	r0, 39
  288=>x"C001",	-- 1100000000000001  li	r1, 0
  289=>x"FFF2",	-- 1111111111110010  liw	r2, font_map + 4 * 0x23
  290=>x"134C",	-- 0001001101001100  
  291=>x"C043",	-- 1100000001000011  li	r3, 8
  292=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  293=>x"01E6",	-- 0000000111100110  
  294=>x"C020",	-- 1100000000100000  li	r0, 4
  295=>x"C001",	-- 1100000000000001  li	r1, 0
  296=>x"FFF2",	-- 1111111111110010  liw	r2, hello_str
  297=>x"16C0",	-- 0001011011000000  
  298=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  299=>x"01A6",	-- 0000000110100110  
  300=>x"2400",	-- 0010010000000000  xor	r0, r0, r0
  301=>x"C0A1",	-- 1100000010100001  li	r1, 20
  302=>x"FFF2",	-- 1111111111110010  liw	r2, 0x2020
  303=>x"2020",	-- 0010000000100000  
  304=>x"D202",	-- 1101001000000010  sw	r2, r0
  305=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  306=>x"FFF2",	-- 1111111111110010  liw	r2, 0x7070
  307=>x"7070",	-- 0111000001110000  
  308=>x"D202",	-- 1101001000000010  sw	r2, r0
  309=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  310=>x"FFF2",	-- 1111111111110010  liw	r2, 0xF8F8
  311=>x"F8F8",	-- 1111100011111000  
  312=>x"D202",	-- 1101001000000010  sw	r2, r0
  313=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  314=>x"FFF2",	-- 1111111111110010  liw	r2, 0xF8F8
  315=>x"F8F8",	-- 1111100011111000  
  316=>x"D202",	-- 1101001000000010  sw	r2, r0
  317=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  318=>x"FFF2",	-- 1111111111110010  liw	r2, 0xF870
  319=>x"F870",	-- 1111100001110000  
  320=>x"D202",	-- 1101001000000010  sw	r2, r0
  321=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  322=>x"FFF2",	-- 1111111111110010  liw	r2, 0x7020
  323=>x"7020",	-- 0111000000100000  
  324=>x"D202",	-- 1101001000000010  sw	r2, r0
  325=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  326=>x"FFF2",	-- 1111111111110010  liw	r2, 0x2070
  327=>x"2070",	-- 0010000001110000  
  328=>x"D202",	-- 1101001000000010  sw	r2, r0
  329=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  330=>x"FFF2",	-- 1111111111110010  liw	r2, 0x0000
  332=>x"D202",	-- 1101001000000010  sw	r2, r0
  333=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  334=>x"C008",	-- 1100000000001000  li	r0, 1
  335=>x"C041",	-- 1100000001000001  li	r1, 8
  336=>x"FFF2",	-- 1111111111110010  liw	r2, font_map
  337=>x"12C0",	-- 0001001011000000  
  338=>x"FFF3",	-- 1111111111110011  liw	r3, PS2_stat
  339=>x"2006",	-- 0010000000000110  
  340=>x"D01B",	-- 1101000000011011  lw	r3, r3
  341=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  342=>x"8824",	-- 1000100000100100  brine	r4, event_not_kbd
  343=>x"063F",	-- 0000011000111111  dec	r7, r7
  344=>x"D23A",	-- 1101001000111010  sw	r2, r7
  345=>x"063F",	-- 0000011000111111  dec	r7, r7
  346=>x"D238",	-- 1101001000111000  sw	r0, r7
  347=>x"063F",	-- 0000011000111111  dec	r7, r7
  348=>x"D239",	-- 1101001000111001  sw	r1, r7
  349=>x"FFF3",	-- 1111111111110011  liw	r3, PS2_rx
  350=>x"2004",	-- 0010000000000100  
  351=>x"D01B",	-- 1101000000011011  lw	r3, r3
  352=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  353=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  354=>x"C043",	-- 1100000001000011  li	r3, 8
  355=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  356=>x"01E6",	-- 0000000111100110  
  357=>x"D039",	-- 1101000000111001  lw	r1, r7
  358=>x"043F",	-- 0000010000111111  inc	r7, r7
  359=>x"D038",	-- 1101000000111000  lw	r0, r7
  360=>x"043F",	-- 0000010000111111  inc	r7, r7
  361=>x"0400",	-- 0000010000000000  inc	r0, r0
  362=>x"C142",	-- 1100000101000010  li	r2, 40
  363=>x"0A82",	-- 0000101010000010  sub	r2, r0, r2
  364=>x"8215",	-- 1000001000010101  brilt	r2, event_kbd_end
  365=>x"6408",	-- 0110010000001000  shr	r0, r1, 2
  366=>x"C042",	-- 1100000001000010  li	r2, 8
  367=>x"0889",	-- 0000100010001001  add	r1, r1, r2
  368=>x"C74A",	-- 1100011101001010  li	r2, 233
  369=>x"0A8A",	-- 0000101010001010  sub	r2, r1, r2
  370=>x"8095",	-- 1000000010010101  brilt	r2, event_kbd_end
  371=>x"C0F1",	-- 1100000011110001  li	r1, 30
  372=>x"D03A",	-- 1101000000111010  lw	r2, r7
  373=>x"043F",	-- 0000010000111111  inc	r7, r7
  374=>x"B703",	-- 1011011100000011  bri	-, event_loop
  375=>x"C750",	-- 1100011101010000  li	r0, 234
  376=>x"C1C2",	-- 1100000111000010  li	r2, 56
  377=>x"FAC6",	-- 1111101011000110  bail	-, r6, div_16_16
  378=>x"018F",	-- 0000000110001111  
  379=>x"C448",	-- 1100010001001000  li	r0, 137
  380=>x"C472",	-- 1100010001110010  li	r2, 142
  381=>x"FAC6",	-- 1111101011000110  bail	-, r6, mult_16_16
  382=>x"0183",	-- 0000000110000011  
  383=>x"C03A",	-- 1100000000111010  li r2, 7
  384=>x"FAC6",	-- 1111101011000110  bail	-, r6, fact_16
  385=>x"019A",	-- 0000000110011010  
  386=>x"FFFF",	-- 1111111111111111  reset
  387=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  388=>x"2524",	-- 0010010100100100  xor	r4, r4, r4
  389=>x"C085",	-- 1100000010000101  li	r5, 16
  390=>x"0849",	-- 0000100001001001  add	r1, r1, r1
  391=>x"0C00",	-- 0000110000000000  adc	r0, r0, r0
  392=>x"0EDB",	-- 0000111011011011  sbc	r3, r3, r3
  393=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  394=>x"08C9",	-- 0000100011001001  add	r1, r1, r3
  395=>x"0D00",	-- 0000110100000000  adc	r0, r0, r4
  396=>x"062D",	-- 0000011000101101  dec	r5, r5
  397=>x"BE6C",	-- 1011111001101100  brine	r5, mult_16_16.loop
  398=>x"E383",	-- 1110001110000011  ba	-, r6
  399=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  400=>x"C084",	-- 1100000010000100  li	r4, 16
  401=>x"0800",	-- 0000100000000000  add	r0, r0, r0
  402=>x"0C49",	-- 0000110001001001  adc	r1, r1, r1
  403=>x"0A8B",	-- 0000101010001011  sub	r3, r1, r2
  404=>x"80DD",	-- 1000000011011101  brilt	r3, div_16_16.skip
  405=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  406=>x"0400",	-- 0000010000000000  inc	r0, r0
  407=>x"0624",	-- 0000011000100100  dec	r4, r4
  408=>x"BE64",	-- 1011111001100100  brine	r4, div_16_16.loop
  409=>x"E383",	-- 1110001110000011  ba	-, r6
  410=>x"2400",	-- 0010010000000000  xor	r0, r0, r0
  411=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  412=>x"8250",	-- 1000001001010000  brieq	r2, fact_16.end
  413=>x"0409",	-- 0000010000001001  inc	r1, r1
  414=>x"1008",	-- 0001000000001000  mova	r0, r1
  415=>x"FAC6",	-- 1111101011000110  bail	-, r6, mult_16_16
  416=>x"0183",	-- 0000000110000011  
  417=>x"8104",	-- 1000000100000100  brine	r0, fact_16.overflow
  418=>x"0183",	-- 0000000110000011  
  419=>x"0612",	-- 0000011000010010  dec	r2, r2
  420=>x"BE94",	-- 1011111010010100  brine	r2, fact_16.loop
  421=>x"E383",	-- 1110001110000011  ba	-, r6
  422=>x"063F",	-- 0000011000111111  dec	r7, r7
  423=>x"D23E",	-- 1101001000111110  sw	r6, r7
  424=>x"D013",	-- 1101000000010011  lw	r3, r2
  425=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  426=>x"8B98",	-- 1000101110011000  brieq	r3, puts.end
  427=>x"063F",	-- 0000011000111111  dec	r7, r7
  428=>x"D238",	-- 1101001000111000  sw	r0, r7
  429=>x"063F",	-- 0000011000111111  dec	r7, r7
  430=>x"D239",	-- 1101001000111001  sw	r1, r7
  431=>x"063F",	-- 0000011000111111  dec	r7, r7
  432=>x"D23A",	-- 1101001000111010  sw	r2, r7
  433=>x"FFF4",	-- 1111111111110100  liw	r4, font_map
  434=>x"12C0",	-- 0001001011000000  
  435=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  436=>x"091A",	-- 0000100100011010  add	r2, r3, r4
  437=>x"C043",	-- 1100000001000011  li	r3, 8
  438=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  439=>x"01E6",	-- 0000000111100110  
  440=>x"D03A",	-- 1101000000111010  lw	r2, r7
  441=>x"043F",	-- 0000010000111111  inc	r7, r7
  442=>x"D039",	-- 1101000000111001  lw	r1, r7
  443=>x"043F",	-- 0000010000111111  inc	r7, r7
  444=>x"D038",	-- 1101000000111000  lw	r0, r7
  445=>x"043F",	-- 0000010000111111  inc	r7, r7
  446=>x"0400",	-- 0000010000000000  inc	r0, r0
  447=>x"D013",	-- 1101000000010011  lw	r3, r2
  448=>x"4E1B",	-- 0100111000011011  shl	r3, r3, 7
  449=>x"6A1B",	-- 0110101000011011  shr	r3, r3, 5
  450=>x"8598",	-- 1000010110011000  brieq	r3, puts.end
  451=>x"063F",	-- 0000011000111111  dec	r7, r7
  452=>x"D238",	-- 1101001000111000  sw	r0, r7
  453=>x"063F",	-- 0000011000111111  dec	r7, r7
  454=>x"D239",	-- 1101001000111001  sw	r1, r7
  455=>x"063F",	-- 0000011000111111  dec	r7, r7
  456=>x"D23A",	-- 1101001000111010  sw	r2, r7
  457=>x"FFF4",	-- 1111111111110100  liw	r4, font_map
  458=>x"12C0",	-- 0001001011000000  
  459=>x"091A",	-- 0000100100011010  add	r2, r3, r4
  460=>x"C043",	-- 1100000001000011  li	r3, 8
  461=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  462=>x"01E6",	-- 0000000111100110  
  463=>x"D03A",	-- 1101000000111010  lw	r2, r7
  464=>x"043F",	-- 0000010000111111  inc	r7, r7
  465=>x"D039",	-- 1101000000111001  lw	r1, r7
  466=>x"043F",	-- 0000010000111111  inc	r7, r7
  467=>x"D038",	-- 1101000000111000  lw	r0, r7
  468=>x"043F",	-- 0000010000111111  inc	r7, r7
  469=>x"0400",	-- 0000010000000000  inc	r0, r0
  470=>x"0412",	-- 0000010000010010  inc	r2, r2
  471=>x"B443",	-- 1011010001000011  bri	-, puts.loop
  472=>x"D03E",	-- 1101000000111110  lw	r6, r7
  473=>x"043F",	-- 0000010000111111  inc	r7, r7
  474=>x"E383",	-- 1110001110000011  ba	-, r6
  475=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  476=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  477=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  478=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  479=>x"D011",	-- 1101000000010001  lw	r1, r2
  480=>x"D221",	-- 1101001000100001  sw	r1, r4
  481=>x"0412",	-- 0000010000010010  inc	r2, r2
  482=>x"0424",	-- 0000010000100100  inc	r4, r4
  483=>x"061B",	-- 0000011000011011  dec	r3, r3
  484=>x"BEDC",	-- 1011111011011100  brine	r3, put_sprite_16_aligned.loop
  485=>x"E383",	-- 1110001110000011  ba	-, r6
  486=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  487=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  488=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  489=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  490=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  491=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  492=>x"C0A5",	-- 1100000010100101  li	r5, 20
  493=>x"8404",	-- 1000010000000100  brine	r0, put_sprite_8_aligned.loop1
  494=>x"D010",	-- 1101000000010000  lw	r0, r2
  495=>x"D021",	-- 1101000000100001  lw	r1, r4
  496=>x"1A41",	-- 0001101001000001  mixhl	r1, r0, r1
  497=>x"D221",	-- 1101001000100001  sw	r1, r4
  498=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  499=>x"061B",	-- 0000011000011011  dec	r3, r3
  500=>x"E398",	-- 1110001110011000  baeq	r3, r6
  501=>x"D021",	-- 1101000000100001  lw	r1, r4
  502=>x"1E41",	-- 0001111001000001  mixll	r1, r0, r1
  503=>x"D221",	-- 1101001000100001  sw	r1, r4
  504=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  505=>x"0412",	-- 0000010000010010  inc	r2, r2
  506=>x"061B",	-- 0000011000011011  dec	r3, r3
  507=>x"E398",	-- 1110001110011000  baeq	r3, r6
  508=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop0
  509=>x"D010",	-- 1101000000010000  lw	r0, r2
  510=>x"D021",	-- 1101000000100001  lw	r1, r4
  511=>x"1809",	-- 0001100000001001  mixhh	r1, r1, r0
  512=>x"D221",	-- 1101001000100001  sw	r1, r4
  513=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  514=>x"061B",	-- 0000011000011011  dec	r3, r3
  515=>x"E398",	-- 1110001110011000  baeq	r3, r6
  516=>x"D021",	-- 1101000000100001  lw	r1, r4
  517=>x"1A09",	-- 0001101000001001  mixhl	r1, r1, r0
  518=>x"D221",	-- 1101001000100001  sw	r1, r4
  519=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  520=>x"0412",	-- 0000010000010010  inc	r2, r2
  521=>x"061B",	-- 0000011000011011  dec	r3, r3
  522=>x"E398",	-- 1110001110011000  baeq	r3, r6
  523=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop1
    others => x"0000"
    );
begin
  process(CLK)
  begin
    if (CLK'event AND CLK='1') then
      D <= m(to_integer(unsigned(AD)));
    end if;
  end process;
end Behavioral;
