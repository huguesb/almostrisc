----------------------------------------------------------------------------------
--
-- File retrieved, on 07/02/2010, from :
-- http://sebastien-viardot.imag.fr/Enseignements/Archi1A2s/sources/ROMPROG.vhd
--
-- Slightly altered to get rid of vendor-specific packages and adjust formatting
-- Now auto-filled by asrom script
--
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROMPROG is
  Port ( AD : in  STD_LOGIC_VECTOR (12 downto 0);
         D : out  STD_LOGIC_VECTOR (15 downto 0);
         CLK : in STD_LOGIC);
end ROMPROG;

architecture Behavioral of ROMPROG is
  constant low_address: natural := 0;
  constant high_address: natural := 8192;
  subtype octet is std_logic_vector( 15 downto 0 );
  type zone_memoire is
    array (natural range low_address to high_address-1) of octet;
  constant m: zone_memoire:= (
    0=>x"FFF7",	-- 1111111111110111  liw	r7, IRQ_mask
    1=>x"2000",	-- 0010000000000000  
    2=>x"F8C0",	-- 1111100011000000  bai	-, os_init
    3=>x"0100",	-- 0000000100000000  
   16=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_ack
   17=>x"2002",	-- 0010000000000010  
   18=>x"D001",	-- 1101000000000001  lw	r1, r0
   19=>x"F54A",	-- 1111010101001010  bspl	r2, r1, 5
   20=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_error
   21=>x"0050",	-- 0000000001010000  
   22=>x"F4CA",	-- 1111010011001010  bspl	r2, r1, 3
   23=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_kbd
   24=>x"0060",	-- 0000000001100000  
   25=>x"F40A",	-- 1111010000001010  bspl	r2, r1, 0
   26=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_tmr
   27=>x"0040",	-- 0000000001000000  
   28=>x"D201",	-- 1101001000000001  sw	r1, r0
   29=>x"FFFE",	-- 1111111111111110  reti
   64=>x"263F",	-- 0010011000111111  not r7, r7
   65=>x"D7C0",	-- 1101011111000000  out	r7
   66=>x"E383",	-- 1110001110000011  ba	-, r6
   80=>x"25FF",	-- 0010010111111111  xor	r7, r7, r7
   81=>x"D7C0",	-- 1101011111000000  out	r7
   82=>x"E383",	-- 1110001110000011  ba	-, r6
   96=>x"FFF2",	-- 1111111111110010  liw	r2, PS2_rx
   97=>x"2004",	-- 0010000000000100  
   98=>x"D012",	-- 1101000000010010  lw	r2, r2
   99=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map + 8
  100=>x"1808",	-- 0001100000001000  
  101=>x"D01B",	-- 1101000000011011  lw	r3, r3
  102=>x"1EBF",	-- 0001111010111111  mixll	r7, r7, r2
  103=>x"C04C",	-- 1100000001001100  li	r4, 9
  104=>x"D227",	-- 1101001000100111  sw	r7, r4
  105=>x"C784",	-- 1100011110000100  li	r4, 0xF0
  106=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  107=>x"96E0",	-- 1001011011100000  brieq	r4, int_kbd.release
  108=>x"C704",	-- 1100011100000100  li	r4, 0xE0
  109=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  110=>x"94A0",	-- 1001010010100000  brieq	r4, int_kbd.extended
  111=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  112=>x"8AA4",	-- 1000101010100100  brine	r4, int_kbd_ext
  113=>x"C31C",	-- 1100001100011100  li	r4, 0x63
  114=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  115=>x"80E4",	-- 1000000011100100  brine	r4, int_kbd_notup
  116=>x"C00D",	-- 1100000000001101  li	r5, 1
  117=>x"8E83",	-- 1000111010000011  bri	-, int_kbd_end
  118=>x"C30C",	-- 1100001100001100  li	r4, 0x61
  119=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  120=>x"80E4",	-- 1000000011100100  brine	r4, int_kbd_notleft
  121=>x"C015",	-- 1100000000010101  li	r5, 2
  122=>x"8D43",	-- 1000110101000011  bri	-, int_kbd_end
  123=>x"C304",	-- 1100001100000100  li	r4, 0x60
  124=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  125=>x"80E4",	-- 1000000011100100  brine	r4, int_kbd_notdown
  126=>x"C025",	-- 1100000000100101  li	r5, 4
  127=>x"8C03",	-- 1000110000000011  bri	-, int_kbd_end
  128=>x"C354",	-- 1100001101010100  li	r4, 0x6A
  129=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  130=>x"80E4",	-- 1000000011100100  brine	r4, int_kbd_notright
  131=>x"C045",	-- 1100000001000101  li	r5, 8
  132=>x"8AC3",	-- 1000101011000011  bri	-, int_kbd_end
  133=>x"C0EC",	-- 1100000011101100  li	r4, 0x1D
  134=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  135=>x"80E4",	-- 1000000011100100  brine	r4, int_kbd_notW
  136=>x"C00D",	-- 1100000000001101  li	r5, 1
  137=>x"8983",	-- 1000100110000011  bri	-, int_kbd_end
  138=>x"C0E4",	-- 1100000011100100  li	r4, 0x1C
  139=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  140=>x"80E4",	-- 1000000011100100  brine	r4, int_kbd_notA
  141=>x"C015",	-- 1100000000010101  li	r5, 2
  142=>x"8843",	-- 1000100001000011  bri	-, int_kbd_end
  143=>x"C0DC",	-- 1100000011011100  li	r4, 0x1B
  144=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  145=>x"80E4",	-- 1000000011100100  brine	r4, int_kbd_notS
  146=>x"C025",	-- 1100000000100101  li	r5, 4
  147=>x"8703",	-- 1000011100000011  bri	-, int_kbd_end
  148=>x"C11C",	-- 1100000100011100  li	r4, 0x23
  149=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  150=>x"80E4",	-- 1000000011100100  brine	r4, int_kbd_notD
  151=>x"C045",	-- 1100000001000101  li	r5, 8
  152=>x"85C3",	-- 1000010111000011  bri	-, int_kbd_end
  153=>x"8883",	-- 1000100010000011  bri	-, int_kbd_done
  154=>x"C3AC",	-- 1100001110101100  li	r4, 0x75
  155=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  156=>x"80E4",	-- 1000000011100100  brine	r4, int_kbd_ext_notup
  157=>x"C00D",	-- 1100000000001101  li	r5, 1
  158=>x"8443",	-- 1000010001000011  bri	-, int_kbd_end
  159=>x"C35C",	-- 1100001101011100  li	r4, 0x6B
  160=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  161=>x"80E4",	-- 1000000011100100  brine	r4, int_kbd_ext_notleft
  162=>x"C015",	-- 1100000000010101  li	r5, 2
  163=>x"8303",	-- 1000001100000011  bri	-, int_kbd_end
  164=>x"C394",	-- 1100001110010100  li	r4, 0x72
  165=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  166=>x"80E4",	-- 1000000011100100  brine	r4, int_kbd_ext_notdown
  167=>x"C025",	-- 1100000000100101  li	r5, 4
  168=>x"81C3",	-- 1000000111000011  bri	-, int_kbd_end
  169=>x"C3A4",	-- 1100001110100100  li	r4, 0x74
  170=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  171=>x"80E4",	-- 1000000011100100  brine	r4, int_kbd_ext_notright
  172=>x"C045",	-- 1100000001000101  li	r5, 8
  173=>x"8083",	-- 1000000010000011  bri	-, int_kbd_end
  174=>x"8343",	-- 1000001101000011  bri	-, int_kbd_done
  175=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  176=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  177=>x"1800",	-- 0001100000000000  
  178=>x"D01A",	-- 1101000000011010  lw	r2, r3
  179=>x"80E4",	-- 1000000011100100  brine	r4, int_kbd_maskout
  180=>x"2352",	-- 0010001101010010  or	r2, r2, r5
  181=>x"80C3",	-- 1000000011000011  bri	-, int_kbd_write
  182=>x"262D",	-- 0010011000101101  not	r5, r5
  183=>x"2152",	-- 0010000101010010  and	r2, r2, r5
  184=>x"D21A",	-- 1101001000011010  sw	r2, r3
  185=>x"C053",	-- 1100000001010011  li	r3, 10
  186=>x"D21A",	-- 1101001000011010  sw	r2, r3
  187=>x"C003",	-- 1100000000000011  li	r3, 0
  188=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  189=>x"1808",	-- 0001100000001000  
  190=>x"D223",	-- 1101001000100011  sw	r3, r4
  191=>x"E383",	-- 1110001110000011  ba	-, r6
  192=>x"C014",	-- 1100000000010100  li	r4, 2
  193=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  194=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  195=>x"1808",	-- 0001100000001000  
  196=>x"D223",	-- 1101001000100011  sw	r3, r4
  197=>x"E383",	-- 1110001110000011  ba	-, r6
  198=>x"C00C",	-- 1100000000001100  li	r4, 1
  199=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  200=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  201=>x"1808",	-- 0001100000001000  
  202=>x"D223",	-- 1101001000100011  sw	r3, r4
  203=>x"E383",	-- 1110001110000011  ba	-, r6
  256=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_mask
  257=>x"2000",	-- 0010000000000000  
  258=>x"C0C9",	-- 1100000011001001  li	r1, 0x19
  259=>x"D201",	-- 1101001000000001  sw	r1, r0
  260=>x"0400",	-- 0000010000000000  inc	r0, r0
  261=>x"CFF9",	-- 1100111111111001  li	r1, -1
  262=>x"D201",	-- 1101001000000001  sw	r1, r0
  263=>x"C03A",	-- 1100000000111010  li	r2, 7
  264=>x"0880",	-- 0000100010000000  add	r0, r0, r2
  265=>x"C0EA",	-- 1100000011101010  li	r2, 0x1D
  266=>x"D202",	-- 1101001000000010  sw	r2, r0
  267=>x"0400",	-- 0000010000000000  inc	r0, r0
  268=>x"C07A",	-- 1100000001111010  li	r2, 15
  269=>x"D202",	-- 1101001000000010  sw	r2, r0
  270=>x"FFF0",	-- 1111111111110000  liw	r0, key_press_map
  271=>x"1800",	-- 0001100000000000  
  272=>x"C001",	-- 1100000000000001  li	r1, 0
  273=>x"D201",	-- 1101001000000001  sw	r1, r0
  274=>x"0400",	-- 0000010000000000  inc	r0, r0
  275=>x"D201",	-- 1101001000000001  sw	r1, r0
  276=>x"0400",	-- 0000010000000000  inc	r0, r0
  277=>x"D201",	-- 1101001000000001  sw	r1, r0
  278=>x"0400",	-- 0000010000000000  inc	r0, r0
  279=>x"D201",	-- 1101001000000001  sw	r1, r0
  280=>x"0400",	-- 0000010000000000  inc	r0, r0
  281=>x"D201",	-- 1101001000000001  sw	r1, r0
  282=>x"0400",	-- 0000010000000000  inc	r0, r0
  283=>x"D201",	-- 1101001000000001  sw	r1, r0
  284=>x"0400",	-- 0000010000000000  inc	r0, r0
  285=>x"D201",	-- 1101001000000001  sw	r1, r0
  286=>x"0400",	-- 0000010000000000  inc	r0, r0
  287=>x"D201",	-- 1101001000000001  sw	r1, r0
  288=>x"0400",	-- 0000010000000000  inc	r0, r0
  289=>x"D201",	-- 1101001000000001  sw	r1, r0
  290=>x"C0F3",	-- 1100000011110011  li	r3, 30
  291=>x"CFFA",	-- 1100111111111010  li	r2, -1
  292=>x"D21A",	-- 1101001000011010  sw	r2, r3
  293=>x"FFF0",	-- 1111111111110000  liw	r0, 0x8421
  294=>x"8421",	-- 1000010000100001  
  295=>x"FFF1",	-- 1111111111110001  liw	r1, 0x1234
  296=>x"1234",	-- 0001001000110100  
  297=>x"D640",	-- 1101011001000000  out	r1
  298=>x"E408",	-- 1110010000001000  exw	r0, r1
  299=>x"E408",	-- 1110010000001000  exw	r0, r1
  300=>x"1842",	-- 0001100001000010  mixhh	r2, r0, r1
  301=>x"1A43",	-- 0001101001000011  mixhl	r3, r0, r1
  302=>x"1C44",	-- 0001110001000100  mixlh	r4, r0, r1
  303=>x"1E45",	-- 0001111001000101  mixll	r5, r0, r1
  304=>x"C01E",	-- 1100000000011110  li	r6, 3
  305=>x"3985",	-- 0011100110000101  rrr	r5, r0, r6
  306=>x"3B8D",	-- 0011101110001101  rrl	r5, r1, r6
  307=>x"3D95",	-- 0011110110010101  rsr	r5, r2, r6
  308=>x"3F9D",	-- 0011111110011101  rsl	r5, r3, r6
  309=>x"FC0E",	-- 1111110000001110  mul	r6, r1, r0
  310=>x"C138",	-- 1100000100111000  li	r0, 39
  311=>x"C001",	-- 1100000000000001  li	r1, 0
  312=>x"FFF2",	-- 1111111111110010  liw	r2, font_map + 4 * 0x23
  313=>x"134C",	-- 0001001101001100  
  314=>x"C043",	-- 1100000001000011  li	r3, 8
  315=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  316=>x"0216",	-- 0000001000010110  
  317=>x"C020",	-- 1100000000100000  li	r0, 4
  318=>x"C001",	-- 1100000000000001  li	r1, 0
  319=>x"FFF2",	-- 1111111111110010  liw	r2, hello_str
  320=>x"16C0",	-- 0001011011000000  
  321=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  322=>x"01DC",	-- 0000000111011100  
  323=>x"2400",	-- 0010010000000000  xor	r0, r0, r0
  324=>x"C0A1",	-- 1100000010100001  li	r1, 20
  325=>x"FFF2",	-- 1111111111110010  liw	r2, 0x2020
  326=>x"2020",	-- 0010000000100000  
  327=>x"D202",	-- 1101001000000010  sw	r2, r0
  328=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  329=>x"FFF2",	-- 1111111111110010  liw	r2, 0x7070
  330=>x"7070",	-- 0111000001110000  
  331=>x"D202",	-- 1101001000000010  sw	r2, r0
  332=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  333=>x"FFF2",	-- 1111111111110010  liw	r2, 0xF8F8
  334=>x"F8F8",	-- 1111100011111000  
  335=>x"D202",	-- 1101001000000010  sw	r2, r0
  336=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  337=>x"FFF2",	-- 1111111111110010  liw	r2, 0xF8F8
  338=>x"F8F8",	-- 1111100011111000  
  339=>x"D202",	-- 1101001000000010  sw	r2, r0
  340=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  341=>x"FFF2",	-- 1111111111110010  liw	r2, 0xF870
  342=>x"F870",	-- 1111100001110000  
  343=>x"D202",	-- 1101001000000010  sw	r2, r0
  344=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  345=>x"FFF2",	-- 1111111111110010  liw	r2, 0x7020
  346=>x"7020",	-- 0111000000100000  
  347=>x"D202",	-- 1101001000000010  sw	r2, r0
  348=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  349=>x"FFF2",	-- 1111111111110010  liw	r2, 0x2070
  350=>x"2070",	-- 0010000001110000  
  351=>x"D202",	-- 1101001000000010  sw	r2, r0
  352=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  353=>x"FFF2",	-- 1111111111110010  liw	r2, 0x0000
  355=>x"D202",	-- 1101001000000010  sw	r2, r0
  356=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  357=>x"C040",	-- 1100000001000000  li	r0, 8
  358=>x"C041",	-- 1100000001000001  li	r1, 8
  359=>x"063F",	-- 0000011000111111  dec	r7, r7
  360=>x"D239",	-- 1101001000111001  sw	r1, r7
  361=>x"063F",	-- 0000011000111111  dec	r7, r7
  362=>x"D238",	-- 1101001000111000  sw	r0, r7
  363=>x"FFF2",	-- 1111111111110010  liw	r2, font_map + 4 * 0x23
  364=>x"134C",	-- 0001001101001100  
  365=>x"C043",	-- 1100000001000011  li	r3, 8
  366=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  367=>x"023C",	-- 0000001000111100  
  368=>x"D038",	-- 1101000000111000  lw	r0, r7
  369=>x"043F",	-- 0000010000111111  inc	r7, r7
  370=>x"D039",	-- 1101000000111001  lw	r1, r7
  371=>x"043F",	-- 0000010000111111  inc	r7, r7
  372=>x"C0A2",	-- 1100000010100010  li	r2, 20
  373=>x"C003",	-- 1100000000000011  li	r3, 0
  374=>x"061B",	-- 0000011000011011  dec	r3, r3
  375=>x"BFDC",	-- 1011111111011100  brine	r3, $-1
  376=>x"0612",	-- 0000011000010010  dec	r2, r2
  377=>x"BF14",	-- 1011111100010100  brine	r2, $-4
  378=>x"FFF2",	-- 1111111111110010  liw	r2, key_press_map
  379=>x"1800",	-- 0001100000000000  
  380=>x"D012",	-- 1101000000010010  lw	r2, r2
  381=>x"8BD0",	-- 1000101111010000  brieq	r2, event_not_kbd
  382=>x"063F",	-- 0000011000111111  dec	r7, r7
  383=>x"D23A",	-- 1101001000111010  sw	r2, r7
  384=>x"063F",	-- 0000011000111111  dec	r7, r7
  385=>x"D239",	-- 1101001000111001  sw	r1, r7
  386=>x"063F",	-- 0000011000111111  dec	r7, r7
  387=>x"D238",	-- 1101001000111000  sw	r0, r7
  388=>x"FFF2",	-- 1111111111110010  liw	r2, font_map
  389=>x"12C0",	-- 0001001011000000  
  390=>x"C043",	-- 1100000001000011  li	r3, 8
  391=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  392=>x"023C",	-- 0000001000111100  
  393=>x"D038",	-- 1101000000111000  lw	r0, r7
  394=>x"043F",	-- 0000010000111111  inc	r7, r7
  395=>x"D039",	-- 1101000000111001  lw	r1, r7
  396=>x"043F",	-- 0000010000111111  inc	r7, r7
  397=>x"D03A",	-- 1101000000111010  lw	r2, r7
  398=>x"043F",	-- 0000010000111111  inc	r7, r7
  399=>x"F413",	-- 1111010000010011  bspl	r3, r2, 0
  400=>x"81D8",	-- 1000000111011000  brieq	r3, event_kbd_no_up
  401=>x"C043",	-- 1100000001000011  li	r3, 8
  402=>x"0ACB",	-- 0000101011001011  sub	r3, r1, r3
  403=>x"809C",	-- 1000000010011100  brine	r3, event_kbd_no_clip_up
  404=>x"C781",	-- 1100011110000001  li	r1, 240
  405=>x"C043",	-- 1100000001000011  li	r3, 8
  406=>x"0AC9",	-- 0000101011001001  sub	r1, r1, r3
  407=>x"F453",	-- 1111010001010011  bspl	r3, r2, 1
  408=>x"8118",	-- 1000000100011000  brieq	r3, event_kbd_no_left
  409=>x"8084",	-- 1000000010000100  brine	r0, event_kbd_no_clip_left
  410=>x"C9C0",	-- 1100100111000000  li	r0, 39*8
  411=>x"0600",	-- 0000011000000000  dec	r0, r0
  412=>x"F493",	-- 1111010010010011  bspl	r3, r2, 2
  413=>x"81D8",	-- 1000000111011000  brieq	r3, event_kbd_no_down
  414=>x"C743",	-- 1100011101000011  li	r3, 232
  415=>x"0ACB",	-- 0000101011001011  sub	r3, r1, r3
  416=>x"809D",	-- 1000000010011101  brilt	r3, event_kbd_no_clip_down
  417=>x"C001",	-- 1100000000000001  li	r1, 0
  418=>x"C043",	-- 1100000001000011  li	r3, 8
  419=>x"08C9",	-- 0000100011001001  add	r1, r1, r3
  420=>x"F4D3",	-- 1111010011010011  bspl	r3, r2, 3
  421=>x"8198",	-- 1000000110011000  brieq	r3, event_kbd_no_right
  422=>x"C9C3",	-- 1100100111000011  li	r3, 39*8
  423=>x"0AC3",	-- 0000101011000011  sub	r3, r0, r3
  424=>x"809D",	-- 1000000010011101  brilt	r3, event_kbd_no_clip_right
  425=>x"CFF8",	-- 1100111111111000  li	r0, -1
  426=>x"0400",	-- 0000010000000000  inc	r0, r0
  427=>x"AF03",	-- 1010111100000011  bri	-, redraw
  428=>x"B383",	-- 1011001110000011  bri	-, event_loop
  429=>x"C750",	-- 1100011101010000  li	r0, 234
  430=>x"C1C2",	-- 1100000111000010  li	r2, 56
  431=>x"FAC6",	-- 1111101011000110  bail	-, r6, div_16_16
  432=>x"01C5",	-- 0000000111000101  
  433=>x"C448",	-- 1100010001001000  li	r0, 137
  434=>x"C472",	-- 1100010001110010  li	r2, 142
  435=>x"FAC6",	-- 1111101011000110  bail	-, r6, mult_16_16
  436=>x"01B9",	-- 0000000110111001  
  437=>x"C03A",	-- 1100000000111010  li r2, 7
  438=>x"FAC6",	-- 1111101011000110  bail	-, r6, fact_16
  439=>x"01D0",	-- 0000000111010000  
  440=>x"FFFF",	-- 1111111111111111  reset
  441=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  442=>x"2524",	-- 0010010100100100  xor	r4, r4, r4
  443=>x"C085",	-- 1100000010000101  li	r5, 16
  444=>x"0849",	-- 0000100001001001  add	r1, r1, r1
  445=>x"0C00",	-- 0000110000000000  adc	r0, r0, r0
  446=>x"0EDB",	-- 0000111011011011  sbc	r3, r3, r3
  447=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  448=>x"08C9",	-- 0000100011001001  add	r1, r1, r3
  449=>x"0D00",	-- 0000110100000000  adc	r0, r0, r4
  450=>x"062D",	-- 0000011000101101  dec	r5, r5
  451=>x"BE6C",	-- 1011111001101100  brine	r5, mult_16_16.loop
  452=>x"E383",	-- 1110001110000011  ba	-, r6
  453=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  454=>x"C084",	-- 1100000010000100  li	r4, 16
  455=>x"0800",	-- 0000100000000000  add	r0, r0, r0
  456=>x"0C49",	-- 0000110001001001  adc	r1, r1, r1
  457=>x"0A8B",	-- 0000101010001011  sub	r3, r1, r2
  458=>x"80DD",	-- 1000000011011101  brilt	r3, div_16_16.skip
  459=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  460=>x"0400",	-- 0000010000000000  inc	r0, r0
  461=>x"0624",	-- 0000011000100100  dec	r4, r4
  462=>x"BE64",	-- 1011111001100100  brine	r4, div_16_16.loop
  463=>x"E383",	-- 1110001110000011  ba	-, r6
  464=>x"2400",	-- 0010010000000000  xor	r0, r0, r0
  465=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  466=>x"8250",	-- 1000001001010000  brieq	r2, fact_16.end
  467=>x"0409",	-- 0000010000001001  inc	r1, r1
  468=>x"1008",	-- 0001000000001000  mova	r0, r1
  469=>x"FAC6",	-- 1111101011000110  bail	-, r6, mult_16_16
  470=>x"01B9",	-- 0000000110111001  
  471=>x"8104",	-- 1000000100000100  brine	r0, fact_16.overflow
  472=>x"01B9",	-- 0000000110111001  
  473=>x"0612",	-- 0000011000010010  dec	r2, r2
  474=>x"BE94",	-- 1011111010010100  brine	r2, fact_16.loop
  475=>x"E383",	-- 1110001110000011  ba	-, r6
  476=>x"063F",	-- 0000011000111111  dec	r7, r7
  477=>x"D23E",	-- 1101001000111110  sw	r6, r7
  478=>x"D013",	-- 1101000000010011  lw	r3, r2
  479=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  480=>x"84D8",	-- 1000010011011000  brieq	r3, puts.end
  481=>x"063F",	-- 0000011000111111  dec	r7, r7
  482=>x"D23A",	-- 1101001000111010  sw	r2, r7
  483=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  484=>x"01F6",	-- 0000000111110110  
  485=>x"D03A",	-- 1101000000111010  lw	r2, r7
  486=>x"043F",	-- 0000010000111111  inc	r7, r7
  487=>x"D013",	-- 1101000000010011  lw	r3, r2
  488=>x"4E1B",	-- 0100111000011011  shl	r3, r3, 7
  489=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  490=>x"8258",	-- 1000001001011000  brieq	r3, puts.end
  491=>x"063F",	-- 0000011000111111  dec	r7, r7
  492=>x"D23A",	-- 1101001000111010  sw	r2, r7
  493=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  494=>x"01F6",	-- 0000000111110110  
  495=>x"D03A",	-- 1101000000111010  lw	r2, r7
  496=>x"043F",	-- 0000010000111111  inc	r7, r7
  497=>x"0412",	-- 0000010000010010  inc	r2, r2
  498=>x"BB03",	-- 1011101100000011  bri	-, puts.loop
  499=>x"D03E",	-- 1101000000111110  lw	r6, r7
  500=>x"043F",	-- 0000010000111111  inc	r7, r7
  501=>x"E383",	-- 1110001110000011  ba	-, r6
  502=>x"063F",	-- 0000011000111111  dec	r7, r7
  503=>x"D23E",	-- 1101001000111110  sw	r6, r7
  504=>x"063F",	-- 0000011000111111  dec	r7, r7
  505=>x"D238",	-- 1101001000111000  sw	r0, r7
  506=>x"063F",	-- 0000011000111111  dec	r7, r7
  507=>x"D239",	-- 1101001000111001  sw	r1, r7
  508=>x"FFF2",	-- 1111111111110010  liw	r2, font_map
  509=>x"12C0",	-- 0001001011000000  
  510=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  511=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  512=>x"C043",	-- 1100000001000011  li	r3, 8
  513=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  514=>x"0216",	-- 0000001000010110  
  515=>x"D039",	-- 1101000000111001  lw	r1, r7
  516=>x"043F",	-- 0000010000111111  inc	r7, r7
  517=>x"D038",	-- 1101000000111000  lw	r0, r7
  518=>x"043F",	-- 0000010000111111  inc	r7, r7
  519=>x"0400",	-- 0000010000000000  inc	r0, r0
  520=>x"D03E",	-- 1101000000111110  lw	r6, r7
  521=>x"043F",	-- 0000010000111111  inc	r7, r7
  522=>x"E383",	-- 1110001110000011  ba	-, r6
  523=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  524=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  525=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  526=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  527=>x"D011",	-- 1101000000010001  lw	r1, r2
  528=>x"D221",	-- 1101001000100001  sw	r1, r4
  529=>x"0412",	-- 0000010000010010  inc	r2, r2
  530=>x"0424",	-- 0000010000100100  inc	r4, r4
  531=>x"061B",	-- 0000011000011011  dec	r3, r3
  532=>x"BEDC",	-- 1011111011011100  brine	r3, put_sprite_16_aligned.loop
  533=>x"E383",	-- 1110001110000011  ba	-, r6
  534=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  535=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  536=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  537=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  538=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  539=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  540=>x"C0A5",	-- 1100000010100101  li	r5, 20
  541=>x"8404",	-- 1000010000000100  brine	r0, put_sprite_8_aligned.loop1
  542=>x"D010",	-- 1101000000010000  lw	r0, r2
  543=>x"D021",	-- 1101000000100001  lw	r1, r4
  544=>x"1A41",	-- 0001101001000001  mixhl	r1, r0, r1
  545=>x"D221",	-- 1101001000100001  sw	r1, r4
  546=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  547=>x"061B",	-- 0000011000011011  dec	r3, r3
  548=>x"E398",	-- 1110001110011000  baeq	r3, r6
  549=>x"D021",	-- 1101000000100001  lw	r1, r4
  550=>x"1E41",	-- 0001111001000001  mixll	r1, r0, r1
  551=>x"D221",	-- 1101001000100001  sw	r1, r4
  552=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  553=>x"0412",	-- 0000010000010010  inc	r2, r2
  554=>x"061B",	-- 0000011000011011  dec	r3, r3
  555=>x"E398",	-- 1110001110011000  baeq	r3, r6
  556=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop0
  557=>x"D010",	-- 1101000000010000  lw	r0, r2
  558=>x"D021",	-- 1101000000100001  lw	r1, r4
  559=>x"1809",	-- 0001100000001001  mixhh	r1, r1, r0
  560=>x"D221",	-- 1101001000100001  sw	r1, r4
  561=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  562=>x"061B",	-- 0000011000011011  dec	r3, r3
  563=>x"E398",	-- 1110001110011000  baeq	r3, r6
  564=>x"D021",	-- 1101000000100001  lw	r1, r4
  565=>x"1A09",	-- 0001101000001001  mixhl	r1, r1, r0
  566=>x"D221",	-- 1101001000100001  sw	r1, r4
  567=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  568=>x"0412",	-- 0000010000010010  inc	r2, r2
  569=>x"061B",	-- 0000011000011011  dec	r3, r3
  570=>x"E398",	-- 1110001110011000  baeq	r3, r6
  571=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop1
  572=>x"C03D",	-- 1100000000111101  li	r5, 7
  573=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  574=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  575=>x"B5E8",	-- 1011010111101000  brieq	r5, put_sprite_8_aligned
  576=>x"062D",	-- 0000011000101101  dec	r5, r5
  577=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  578=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  579=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  580=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  581=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  582=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  583=>x"8AC4",	-- 1000101011000100  brine	r0, put_sprite_8.loop1
  584=>x"D010",	-- 1101000000010000  lw	r0, r2
  585=>x"063F",	-- 0000011000111111  dec	r7, r7
  586=>x"D23A",	-- 1101001000111010  sw	r2, r7
  587=>x"C002",	-- 1100000000000010  li	r2, 0
  588=>x"1A80",	-- 0001101010000000  mixhl	r0, r0, r2
  589=>x"C802",	-- 1100100000000010  li	r2, 0x100
  590=>x"3B52",	-- 0011101101010010  rrl	r2, r2, r5
  591=>x"3B40",	-- 0011101101000000  rrl	r0, r0, r5
  592=>x"D021",	-- 1101000000100001  lw	r1, r4
  593=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  594=>x"2612",	-- 0010011000010010  not	r2, r2
  595=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  596=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  597=>x"D221",	-- 1101001000100001  sw	r1, r4
  598=>x"C0A1",	-- 1100000010100001  li	r1, 20
  599=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  600=>x"D03A",	-- 1101000000111010  lw	r2, r7
  601=>x"043F",	-- 0000010000111111  inc	r7, r7
  602=>x"061B",	-- 0000011000011011  dec	r3, r3
  603=>x"E398",	-- 1110001110011000  baeq	r3, r6
  604=>x"D010",	-- 1101000000010000  lw	r0, r2
  605=>x"063F",	-- 0000011000111111  dec	r7, r7
  606=>x"D23A",	-- 1101001000111010  sw	r2, r7
  607=>x"C002",	-- 1100000000000010  li	r2, 0
  608=>x"1E80",	-- 0001111010000000  mixll	r0, r0, r2
  609=>x"C802",	-- 1100100000000010  li	r2, 0x100
  610=>x"3B52",	-- 0011101101010010  rrl	r2, r2, r5
  611=>x"3B43",	-- 0011101101000011  rrl	r3, r0, r5
  612=>x"D021",	-- 1101000000100001  lw	r1, r4
  613=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  614=>x"2612",	-- 0010011000010010  not	r2, r2
  615=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  616=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  617=>x"D221",	-- 1101001000100001  sw	r1, r4
  618=>x"C0A1",	-- 1100000010100001  li	r1, 20
  619=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  620=>x"D03A",	-- 1101000000111010  lw	r2, r7
  621=>x"043F",	-- 0000010000111111  inc	r7, r7
  622=>x"0412",	-- 0000010000010010  inc	r2, r2
  623=>x"061B",	-- 0000011000011011  dec	r3, r3
  624=>x"E398",	-- 1110001110011000  baeq	r3, r6
  625=>x"B5C3",	-- 1011010111000011  bri	-, put_sprite_8.loop0
  626=>x"D010",	-- 1101000000010000  lw	r0, r2
  627=>x"063F",	-- 0000011000111111  dec	r7, r7
  628=>x"D23A",	-- 1101001000111010  sw	r2, r7
  629=>x"063F",	-- 0000011000111111  dec	r7, r7
  630=>x"D23B",	-- 1101001000111011  sw	r3, r7
  631=>x"C002",	-- 1100000000000010  li	r2, 0
  632=>x"1C13",	-- 0001110000010011  mixlh	r3, r2, r0
  633=>x"C7FA",	-- 1100011111111010  li	r2, 0xFF
  634=>x"3F52",	-- 0011111101010010  rsl	r2, r2, r5
  635=>x"3F5B",	-- 0011111101011011  rsl	r3, r3, r5
  636=>x"D021",	-- 1101000000100001  lw	r1, r4
  637=>x"20D3",	-- 0010000011010011  and	r3, r2, r3
  638=>x"2612",	-- 0010011000010010  not	r2, r2
  639=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  640=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  641=>x"D221",	-- 1101001000100001  sw	r1, r4
  642=>x"0424",	-- 0000010000100100  inc	r4, r4
  643=>x"C002",	-- 1100000000000010  li	r2, 0
  644=>x"1A83",	-- 0001101010000011  mixhl	r3, r0, r2
  645=>x"CFFA",	-- 1100111111111010  li	r2, -1
  646=>x"3F52",	-- 0011111101010010  rsl	r2, r2, r5
  647=>x"3F5B",	-- 0011111101011011  rsl	r3, r3, r5
  648=>x"D021",	-- 1101000000100001  lw	r1, r4
  649=>x"20D3",	-- 0010000011010011  and	r3, r2, r3
  650=>x"2612",	-- 0010011000010010  not	r2, r2
  651=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  652=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  653=>x"D221",	-- 1101001000100001  sw	r1, r4
  654=>x"C099",	-- 1100000010011001  li	r1, 19
  655=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  656=>x"D03B",	-- 1101000000111011  lw	r3, r7
  657=>x"043F",	-- 0000010000111111  inc	r7, r7
  658=>x"D03A",	-- 1101000000111010  lw	r2, r7
  659=>x"043F",	-- 0000010000111111  inc	r7, r7
  660=>x"061B",	-- 0000011000011011  dec	r3, r3
  661=>x"E398",	-- 1110001110011000  baeq	r3, r6
  662=>x"063F",	-- 0000011000111111  dec	r7, r7
  663=>x"D23A",	-- 1101001000111010  sw	r2, r7
  664=>x"063F",	-- 0000011000111111  dec	r7, r7
  665=>x"D23B",	-- 1101001000111011  sw	r3, r7
  666=>x"C002",	-- 1100000000000010  li	r2, 0
  667=>x"1E13",	-- 0001111000010011  mixll	r3, r2, r0
  668=>x"C7FA",	-- 1100011111111010  li	r2, 0xFF
  669=>x"3F52",	-- 0011111101010010  rsl	r2, r2, r5
  670=>x"3F5B",	-- 0011111101011011  rsl	r3, r3, r5
  671=>x"D021",	-- 1101000000100001  lw	r1, r4
  672=>x"20D3",	-- 0010000011010011  and	r3, r2, r3
  673=>x"2612",	-- 0010011000010010  not	r2, r2
  674=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  675=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  676=>x"D221",	-- 1101001000100001  sw	r1, r4
  677=>x"0424",	-- 0000010000100100  inc	r4, r4
  678=>x"C002",	-- 1100000000000010  li	r2, 0
  679=>x"1E83",	-- 0001111010000011  mixll	r3, r0, r2
  680=>x"CFFA",	-- 1100111111111010  li	r2, -1
  681=>x"3F52",	-- 0011111101010010  rsl	r2, r2, r5
  682=>x"3F5B",	-- 0011111101011011  rsl	r3, r3, r5
  683=>x"D021",	-- 1101000000100001  lw	r1, r4
  684=>x"20D3",	-- 0010000011010011  and	r3, r2, r3
  685=>x"2612",	-- 0010011000010010  not	r2, r2
  686=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  687=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  688=>x"D221",	-- 1101001000100001  sw	r1, r4
  689=>x"C0E9",	-- 1100000011101001  li	r1, 29
  690=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  691=>x"D03B",	-- 1101000000111011  lw	r3, r7
  692=>x"043F",	-- 0000010000111111  inc	r7, r7
  693=>x"D03A",	-- 1101000000111010  lw	r2, r7
  694=>x"043F",	-- 0000010000111111  inc	r7, r7
  695=>x"0412",	-- 0000010000010010  inc	r2, r2
  696=>x"061B",	-- 0000011000011011  dec	r3, r3
  697=>x"E398",	-- 1110001110011000  baeq	r3, r6
  698=>x"AE03",	-- 1010111000000011  bri	-, put_sprite_8.loop1
    others => x"0000"
    );
begin
  process(CLK)
  begin
    if (CLK'event AND CLK='1') then
      D <= m(to_integer(unsigned(AD)));
    end if;
  end process;
end Behavioral;
