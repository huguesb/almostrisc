----------------------------------------------------------------------------------
--
-- File retrieved, on 07/02/2010, from :
-- http://sebastien-viardot.imag.fr/Enseignements/Archi1A2s/sources/RAMDoublePort.vhd
--
-- Slightly altered to get rid of vendor-specific packages and adjust formatting
-- Now auto-filled by asrom script
--
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity RAMDoublePort is
    Port ( AD1 : in  STD_LOGIC_VECTOR (12 downto 0);
           AD2 : in  STD_LOGIC_VECTOR (12 downto 0);
           DIN1 : in  STD_LOGIC_VECTOR (15 downto 0);
           DOUT1 : out  STD_LOGIC_VECTOR (15 downto 0);
           WE1 : in  STD_LOGIC;
           DOUT2 : out  STD_LOGIC_VECTOR (15 downto 0);
           OE1 : in  STD_LOGIC;
           CE1 : in  STD_LOGIC;
			  CLK : in STD_LOGIC);
end RAMDoublePort;

 -- memory map :
 --     0 -  4799 : VGA-mapped RAM (320*240 pix, 16 pix per word => 4800 words)
 --  4800 -  5823 : font map (8*8 : 4 words per character, 256 chars => 1024 words)
 --  5824 -  8191 : user data (2368 words)

architecture Behavioral of RAMDoublePort is
 constant low_address: natural := 0;
 constant high_address: natural := 8192;  
 subtype octet is std_logic_vector( 15 downto 0 );
 type zone_memoire is
         array (natural range low_address to high_address) of octet;
 signal memoire: zone_memoire := (
     0 => x"0000",
     1 => x"0000",
     2 => x"0000",
     3 => x"0000",
     4 => x"0000",
     5 => x"0000",
     6 => x"0000",
     7 => x"0000",
     8 => x"0000",
     9 => x"0000",
    10 => x"0000",
    11 => x"0000",
    12 => x"0000",
    13 => x"0000",
    14 => x"0000",
    15 => x"0000",
    16 => x"0000",
    17 => x"0000",
    18 => x"0000",
    19 => x"0000",
    20 => x"0000",
    21 => x"0000",
    22 => x"0000",
    23 => x"0000",
    24 => x"0000",
    25 => x"0000",
    26 => x"0000",
    27 => x"0000",
    28 => x"0000",
    29 => x"0000",
    30 => x"0000",
    31 => x"0000",
    32 => x"0000",
    33 => x"0000",
    34 => x"0000",
    35 => x"0000",
    36 => x"0000",
    37 => x"0000",
    38 => x"0000",
    39 => x"0000",
    40 => x"0000",
    41 => x"0000",
    42 => x"0000",
    43 => x"0000",
    44 => x"0000",
    45 => x"0000",
    46 => x"0000",
    47 => x"0000",
    48 => x"0000",
    49 => x"0000",
    50 => x"0000",
    51 => x"0000",
    52 => x"0000",
    53 => x"0000",
    54 => x"0000",
    55 => x"0000",
    56 => x"0000",
    57 => x"0000",
    58 => x"0000",
    59 => x"0000",
    60 => x"0000",
    61 => x"0000",
    62 => x"0000",
    63 => x"0000",
    64 => x"0000",
    65 => x"0000",
    66 => x"0000",
    67 => x"0000",
    68 => x"0000",
    69 => x"0000",
    70 => x"0000",
    71 => x"0000",
    72 => x"0000",
    73 => x"0000",
    74 => x"0000",
    75 => x"0000",
    76 => x"0000",
    77 => x"0000",
    78 => x"0000",
    79 => x"0000",
    80 => x"0000",
    81 => x"0000",
    82 => x"0000",
    83 => x"0000",
    84 => x"0000",
    85 => x"0000",
    86 => x"0000",
    87 => x"0000",
    88 => x"0000",
    89 => x"0000",
    90 => x"0000",
    91 => x"0000",
    92 => x"0000",
    93 => x"0000",
    94 => x"0000",
    95 => x"0000",
    96 => x"0000",
    97 => x"0000",
    98 => x"0000",
    99 => x"0000",
   100 => x"0000",
   101 => x"0000",
   102 => x"0000",
   103 => x"0000",
   104 => x"0000",
   105 => x"0000",
   106 => x"0000",
   107 => x"0000",
   108 => x"0000",
   109 => x"0000",
   110 => x"0000",
   111 => x"0000",
   112 => x"0000",
   113 => x"0000",
   114 => x"0000",
   115 => x"0000",
   116 => x"0000",
   117 => x"0000",
   118 => x"0000",
   119 => x"0000",
   120 => x"0000",
   121 => x"0000",
   122 => x"0000",
   123 => x"0000",
   124 => x"0000",
   125 => x"0000",
   126 => x"0000",
   127 => x"0000",
   128 => x"0000",
   129 => x"0000",
   130 => x"0000",
   131 => x"0000",
   132 => x"0000",
   133 => x"0000",
   134 => x"0000",
   135 => x"0000",
   136 => x"0000",
   137 => x"0000",
   138 => x"0000",
   139 => x"0000",
   140 => x"0000",
   141 => x"0000",
   142 => x"0000",
   143 => x"0000",
   144 => x"0000",
   145 => x"0000",
   146 => x"0000",
   147 => x"0000",
   148 => x"0000",
   149 => x"0000",
   150 => x"0000",
   151 => x"0000",
   152 => x"0000",
   153 => x"0000",
   154 => x"0000",
   155 => x"0000",
   156 => x"0000",
   157 => x"0000",
   158 => x"0000",
   159 => x"0000",
   160 => x"0000",
   161 => x"0000",
   162 => x"0000",
   163 => x"0000",
   164 => x"0000",
   165 => x"0000",
   166 => x"0000",
   167 => x"0000",
   168 => x"0000",
   169 => x"0000",
   170 => x"0000",
   171 => x"0000",
   172 => x"0000",
   173 => x"0000",
   174 => x"0000",
   175 => x"0000",
   176 => x"0000",
   177 => x"0000",
   178 => x"0000",
   179 => x"0000",
   180 => x"0000",
   181 => x"0000",
   182 => x"0000",
   183 => x"0000",
   184 => x"0000",
   185 => x"0000",
   186 => x"0000",
   187 => x"0000",
   188 => x"0000",
   189 => x"0000",
   190 => x"0000",
   191 => x"0000",
   192 => x"0000",
   193 => x"0000",
   194 => x"0000",
   195 => x"0000",
   196 => x"0000",
   197 => x"0000",
   198 => x"0000",
   199 => x"0000",
   200 => x"0000",
   201 => x"0000",
   202 => x"0000",
   203 => x"0000",
   204 => x"0000",
   205 => x"0000",
   206 => x"0000",
   207 => x"0000",
   208 => x"0000",
   209 => x"0000",
   210 => x"0000",
   211 => x"0000",
   212 => x"0000",
   213 => x"0000",
   214 => x"0000",
   215 => x"0000",
   216 => x"0000",
   217 => x"0000",
   218 => x"0000",
   219 => x"0000",
   220 => x"0000",
   221 => x"0000",
   222 => x"0000",
   223 => x"0000",
   224 => x"0000",
   225 => x"0000",
   226 => x"0000",
   227 => x"0000",
   228 => x"0000",
   229 => x"0000",
   230 => x"0000",
   231 => x"0000",
   232 => x"0000",
   233 => x"0000",
   234 => x"0000",
   235 => x"0000",
   236 => x"0000",
   237 => x"0000",
   238 => x"0000",
   239 => x"0000",
   240 => x"0000",
   241 => x"0000",
   242 => x"0000",
   243 => x"0000",
   244 => x"0000",
   245 => x"0000",
   246 => x"0000",
   247 => x"0000",
   248 => x"0000",
   249 => x"0000",
   250 => x"0000",
   251 => x"0000",
   252 => x"0000",
   253 => x"0000",
   254 => x"0000",
   255 => x"0000",
   256 => x"0000",
   257 => x"0000",
   258 => x"0000",
   259 => x"0000",
   260 => x"0000",
   261 => x"0000",
   262 => x"0000",
   263 => x"0000",
   264 => x"0000",
   265 => x"0000",
   266 => x"0000",
   267 => x"0000",
   268 => x"0000",
   269 => x"0000",
   270 => x"0000",
   271 => x"0000",
   272 => x"0000",
   273 => x"0000",
   274 => x"0000",
   275 => x"0000",
   276 => x"0000",
   277 => x"0000",
   278 => x"0000",
   279 => x"0000",
   280 => x"0000",
   281 => x"0000",
   282 => x"0000",
   283 => x"0000",
   284 => x"0000",
   285 => x"0000",
   286 => x"0000",
   287 => x"0000",
   288 => x"0000",
   289 => x"0000",
   290 => x"0000",
   291 => x"0000",
   292 => x"0000",
   293 => x"0000",
   294 => x"0000",
   295 => x"0000",
   296 => x"0000",
   297 => x"0000",
   298 => x"0000",
   299 => x"0000",
   300 => x"0000",
   301 => x"0000",
   302 => x"0000",
   303 => x"0000",
   304 => x"0000",
   305 => x"0000",
   306 => x"0000",
   307 => x"0000",
   308 => x"0000",
   309 => x"0000",
   310 => x"0000",
   311 => x"0000",
   312 => x"0000",
   313 => x"0000",
   314 => x"0000",
   315 => x"0000",
   316 => x"0000",
   317 => x"0000",
   318 => x"0000",
   319 => x"0000",
   320 => x"0000",
   321 => x"0000",
   322 => x"0000",
   323 => x"0000",
   324 => x"0000",
   325 => x"0000",
   326 => x"0000",
   327 => x"0000",
   328 => x"0000",
   329 => x"0000",
   330 => x"0000",
   331 => x"0000",
   332 => x"0000",
   333 => x"0000",
   334 => x"0000",
   335 => x"0000",
   336 => x"0000",
   337 => x"0000",
   338 => x"0000",
   339 => x"0000",
   340 => x"0000",
   341 => x"0000",
   342 => x"0000",
   343 => x"0000",
   344 => x"0000",
   345 => x"0000",
   346 => x"0000",
   347 => x"0000",
   348 => x"0000",
   349 => x"0000",
   350 => x"0000",
   351 => x"0000",
   352 => x"0000",
   353 => x"0000",
   354 => x"0000",
   355 => x"0000",
   356 => x"0000",
   357 => x"0000",
   358 => x"0000",
   359 => x"0000",
   360 => x"0000",
   361 => x"0000",
   362 => x"0000",
   363 => x"0000",
   364 => x"0000",
   365 => x"0000",
   366 => x"0000",
   367 => x"0000",
   368 => x"0000",
   369 => x"0000",
   370 => x"0000",
   371 => x"0000",
   372 => x"0000",
   373 => x"0000",
   374 => x"0000",
   375 => x"0000",
   376 => x"0000",
   377 => x"0000",
   378 => x"0000",
   379 => x"0000",
   380 => x"0000",
   381 => x"0000",
   382 => x"0000",
   383 => x"0000",
   384 => x"0000",
   385 => x"0000",
   386 => x"0000",
   387 => x"0000",
   388 => x"0000",
   389 => x"0000",
   390 => x"0000",
   391 => x"0000",
   392 => x"0000",
   393 => x"0000",
   394 => x"0000",
   395 => x"0000",
   396 => x"0000",
   397 => x"0000",
   398 => x"0000",
   399 => x"0000",
   400 => x"0000",
   401 => x"0000",
   402 => x"0000",
   403 => x"0000",
   404 => x"0000",
   405 => x"0000",
   406 => x"0000",
   407 => x"0000",
   408 => x"0000",
   409 => x"0000",
   410 => x"0000",
   411 => x"0000",
   412 => x"0000",
   413 => x"0000",
   414 => x"0000",
   415 => x"0000",
   416 => x"0000",
   417 => x"0000",
   418 => x"0000",
   419 => x"0000",
   420 => x"0000",
   421 => x"0000",
   422 => x"0000",
   423 => x"0000",
   424 => x"0000",
   425 => x"0000",
   426 => x"0000",
   427 => x"0000",
   428 => x"0000",
   429 => x"0000",
   430 => x"0000",
   431 => x"0000",
   432 => x"0000",
   433 => x"0000",
   434 => x"0000",
   435 => x"0000",
   436 => x"0000",
   437 => x"0000",
   438 => x"0000",
   439 => x"0000",
   440 => x"0000",
   441 => x"0000",
   442 => x"0000",
   443 => x"0000",
   444 => x"0000",
   445 => x"0000",
   446 => x"0000",
   447 => x"0000",
   448 => x"0000",
   449 => x"0000",
   450 => x"0000",
   451 => x"0000",
   452 => x"0000",
   453 => x"0000",
   454 => x"0000",
   455 => x"0000",
   456 => x"0000",
   457 => x"0000",
   458 => x"0000",
   459 => x"0000",
   460 => x"0000",
   461 => x"0000",
   462 => x"0000",
   463 => x"0000",
   464 => x"0000",
   465 => x"0000",
   466 => x"0000",
   467 => x"0000",
   468 => x"0000",
   469 => x"0000",
   470 => x"0000",
   471 => x"0000",
   472 => x"0000",
   473 => x"0000",
   474 => x"0000",
   475 => x"0000",
   476 => x"0000",
   477 => x"0000",
   478 => x"0000",
   479 => x"0000",
   480 => x"0000",
   481 => x"0000",
   482 => x"0000",
   483 => x"0000",
   484 => x"0000",
   485 => x"0000",
   486 => x"0000",
   487 => x"0000",
   488 => x"0000",
   489 => x"0000",
   490 => x"0000",
   491 => x"0000",
   492 => x"0000",
   493 => x"0000",
   494 => x"0000",
   495 => x"0000",
   496 => x"0000",
   497 => x"0000",
   498 => x"0000",
   499 => x"0000",
   500 => x"0000",
   501 => x"0000",
   502 => x"0000",
   503 => x"0000",
   504 => x"0000",
   505 => x"0000",
   506 => x"0000",
   507 => x"0000",
   508 => x"0000",
   509 => x"0000",
   510 => x"0000",
   511 => x"0000",
   512 => x"0000",
   513 => x"0000",
   514 => x"0000",
   515 => x"0000",
   516 => x"0000",
   517 => x"0000",
   518 => x"0000",
   519 => x"0000",
   520 => x"0000",
   521 => x"0000",
   522 => x"0000",
   523 => x"0000",
   524 => x"0000",
   525 => x"0000",
   526 => x"0000",
   527 => x"0000",
   528 => x"0000",
   529 => x"0000",
   530 => x"0000",
   531 => x"0000",
   532 => x"0000",
   533 => x"0000",
   534 => x"0000",
   535 => x"0000",
   536 => x"0000",
   537 => x"0000",
   538 => x"0000",
   539 => x"0000",
   540 => x"0000",
   541 => x"0000",
   542 => x"0000",
   543 => x"0000",
   544 => x"0000",
   545 => x"0000",
   546 => x"0000",
   547 => x"0000",
   548 => x"0000",
   549 => x"0000",
   550 => x"0000",
   551 => x"0000",
   552 => x"0000",
   553 => x"0000",
   554 => x"0000",
   555 => x"0000",
   556 => x"0000",
   557 => x"0000",
   558 => x"0000",
   559 => x"0000",
   560 => x"0000",
   561 => x"0000",
   562 => x"0000",
   563 => x"0000",
   564 => x"0000",
   565 => x"0000",
   566 => x"0000",
   567 => x"0000",
   568 => x"0000",
   569 => x"0000",
   570 => x"0000",
   571 => x"0000",
   572 => x"0000",
   573 => x"0000",
   574 => x"0000",
   575 => x"0000",
   576 => x"0000",
   577 => x"0000",
   578 => x"0000",
   579 => x"0000",
   580 => x"0000",
   581 => x"0000",
   582 => x"0000",
   583 => x"0000",
   584 => x"0000",
   585 => x"0000",
   586 => x"0000",
   587 => x"0000",
   588 => x"0000",
   589 => x"0000",
   590 => x"0000",
   591 => x"0000",
   592 => x"0000",
   593 => x"0000",
   594 => x"0000",
   595 => x"0000",
   596 => x"0000",
   597 => x"0000",
   598 => x"0000",
   599 => x"0000",
   600 => x"0000",
   601 => x"0000",
   602 => x"0000",
   603 => x"0000",
   604 => x"0000",
   605 => x"0000",
   606 => x"0000",
   607 => x"0000",
   608 => x"0000",
   609 => x"0000",
   610 => x"0000",
   611 => x"0000",
   612 => x"0000",
   613 => x"0000",
   614 => x"0000",
   615 => x"0000",
   616 => x"0000",
   617 => x"0000",
   618 => x"0000",
   619 => x"0000",
   620 => x"0000",
   621 => x"0000",
   622 => x"0000",
   623 => x"0000",
   624 => x"0000",
   625 => x"0000",
   626 => x"0000",
   627 => x"0000",
   628 => x"0000",
   629 => x"0000",
   630 => x"0000",
   631 => x"0000",
   632 => x"0000",
   633 => x"0000",
   634 => x"0000",
   635 => x"0000",
   636 => x"0000",
   637 => x"0000",
   638 => x"0000",
   639 => x"0000",
   640 => x"0000",
   641 => x"0000",
   642 => x"0000",
   643 => x"0000",
   644 => x"0000",
   645 => x"0000",
   646 => x"0000",
   647 => x"0000",
   648 => x"0000",
   649 => x"0000",
   650 => x"0000",
   651 => x"0000",
   652 => x"0000",
   653 => x"0000",
   654 => x"0000",
   655 => x"0000",
   656 => x"0000",
   657 => x"0000",
   658 => x"0000",
   659 => x"0000",
   660 => x"0000",
   661 => x"0000",
   662 => x"0000",
   663 => x"0000",
   664 => x"0000",
   665 => x"0000",
   666 => x"0000",
   667 => x"0000",
   668 => x"0000",
   669 => x"0000",
   670 => x"0000",
   671 => x"0000",
   672 => x"0000",
   673 => x"0000",
   674 => x"0000",
   675 => x"0000",
   676 => x"0000",
   677 => x"0000",
   678 => x"0000",
   679 => x"0000",
   680 => x"0000",
   681 => x"0000",
   682 => x"0000",
   683 => x"0000",
   684 => x"0000",
   685 => x"0000",
   686 => x"0000",
   687 => x"0000",
   688 => x"0000",
   689 => x"0000",
   690 => x"0000",
   691 => x"0000",
   692 => x"0000",
   693 => x"0000",
   694 => x"0000",
   695 => x"0000",
   696 => x"0000",
   697 => x"0000",
   698 => x"0000",
   699 => x"0000",
   700 => x"0000",
   701 => x"0000",
   702 => x"0000",
   703 => x"0000",
   704 => x"0000",
   705 => x"0000",
   706 => x"0000",
   707 => x"0000",
   708 => x"0000",
   709 => x"0000",
   710 => x"0000",
   711 => x"0000",
   712 => x"0000",
   713 => x"0000",
   714 => x"0000",
   715 => x"0000",
   716 => x"0000",
   717 => x"0000",
   718 => x"0000",
   719 => x"0000",
   720 => x"0000",
   721 => x"0000",
   722 => x"0000",
   723 => x"0000",
   724 => x"0000",
   725 => x"0000",
   726 => x"0000",
   727 => x"0000",
   728 => x"0000",
   729 => x"0000",
   730 => x"0000",
   731 => x"0000",
   732 => x"0000",
   733 => x"0000",
   734 => x"0000",
   735 => x"0000",
   736 => x"0000",
   737 => x"0000",
   738 => x"0000",
   739 => x"0000",
   740 => x"0000",
   741 => x"0000",
   742 => x"0000",
   743 => x"0000",
   744 => x"0000",
   745 => x"0000",
   746 => x"0000",
   747 => x"0000",
   748 => x"0000",
   749 => x"0000",
   750 => x"0000",
   751 => x"0000",
   752 => x"0000",
   753 => x"0000",
   754 => x"0000",
   755 => x"0000",
   756 => x"0000",
   757 => x"0000",
   758 => x"0000",
   759 => x"0000",
   760 => x"0000",
   761 => x"0000",
   762 => x"0000",
   763 => x"0000",
   764 => x"0000",
   765 => x"0000",
   766 => x"0000",
   767 => x"0000",
   768 => x"0000",
   769 => x"0000",
   770 => x"0000",
   771 => x"0000",
   772 => x"0000",
   773 => x"0000",
   774 => x"0000",
   775 => x"0000",
   776 => x"0000",
   777 => x"0000",
   778 => x"0000",
   779 => x"0000",
   780 => x"0000",
   781 => x"0000",
   782 => x"0000",
   783 => x"0000",
   784 => x"0000",
   785 => x"0000",
   786 => x"0000",
   787 => x"0000",
   788 => x"0000",
   789 => x"0000",
   790 => x"0000",
   791 => x"0000",
   792 => x"0000",
   793 => x"0000",
   794 => x"0000",
   795 => x"0000",
   796 => x"0000",
   797 => x"0000",
   798 => x"0000",
   799 => x"0000",
   800 => x"0000",
   801 => x"0000",
   802 => x"0000",
   803 => x"0000",
   804 => x"0000",
   805 => x"0000",
   806 => x"0000",
   807 => x"0000",
   808 => x"0000",
   809 => x"0000",
   810 => x"0000",
   811 => x"0000",
   812 => x"0000",
   813 => x"0000",
   814 => x"0000",
   815 => x"0000",
   816 => x"0000",
   817 => x"0000",
   818 => x"0000",
   819 => x"0000",
   820 => x"0000",
   821 => x"0000",
   822 => x"0000",
   823 => x"0000",
   824 => x"0000",
   825 => x"0000",
   826 => x"0000",
   827 => x"0000",
   828 => x"0000",
   829 => x"0000",
   830 => x"0000",
   831 => x"0000",
   832 => x"0000",
   833 => x"0000",
   834 => x"0000",
   835 => x"0000",
   836 => x"0000",
   837 => x"0000",
   838 => x"0000",
   839 => x"0000",
   840 => x"0000",
   841 => x"0000",
   842 => x"0000",
   843 => x"0000",
   844 => x"0000",
   845 => x"0000",
   846 => x"0000",
   847 => x"0000",
   848 => x"0000",
   849 => x"0000",
   850 => x"0000",
   851 => x"0000",
   852 => x"0000",
   853 => x"0000",
   854 => x"0000",
   855 => x"0000",
   856 => x"0000",
   857 => x"0000",
   858 => x"0000",
   859 => x"0000",
   860 => x"0000",
   861 => x"0000",
   862 => x"0000",
   863 => x"0000",
   864 => x"0000",
   865 => x"0000",
   866 => x"0000",
   867 => x"0000",
   868 => x"0000",
   869 => x"0000",
   870 => x"0000",
   871 => x"0000",
   872 => x"0000",
   873 => x"0000",
   874 => x"0000",
   875 => x"0000",
   876 => x"0000",
   877 => x"0000",
   878 => x"0000",
   879 => x"0000",
   880 => x"0000",
   881 => x"0000",
   882 => x"0000",
   883 => x"0000",
   884 => x"0000",
   885 => x"0000",
   886 => x"0000",
   887 => x"0000",
   888 => x"0000",
   889 => x"0000",
   890 => x"0000",
   891 => x"0000",
   892 => x"0000",
   893 => x"0000",
   894 => x"0000",
   895 => x"0000",
   896 => x"0000",
   897 => x"0000",
   898 => x"0000",
   899 => x"0000",
   900 => x"0000",
   901 => x"0000",
   902 => x"0000",
   903 => x"0000",
   904 => x"0000",
   905 => x"0000",
   906 => x"0000",
   907 => x"0000",
   908 => x"0000",
   909 => x"0000",
   910 => x"0000",
   911 => x"0000",
   912 => x"0000",
   913 => x"0000",
   914 => x"0000",
   915 => x"0000",
   916 => x"0000",
   917 => x"0000",
   918 => x"0000",
   919 => x"0000",
   920 => x"0000",
   921 => x"0000",
   922 => x"0000",
   923 => x"0000",
   924 => x"0000",
   925 => x"0000",
   926 => x"0000",
   927 => x"0000",
   928 => x"0000",
   929 => x"0000",
   930 => x"0000",
   931 => x"0000",
   932 => x"0000",
   933 => x"0000",
   934 => x"0000",
   935 => x"0000",
   936 => x"0000",
   937 => x"0000",
   938 => x"0000",
   939 => x"0000",
   940 => x"0000",
   941 => x"0000",
   942 => x"0000",
   943 => x"0000",
   944 => x"0000",
   945 => x"0000",
   946 => x"0000",
   947 => x"0000",
   948 => x"0000",
   949 => x"0000",
   950 => x"0000",
   951 => x"0000",
   952 => x"0000",
   953 => x"0000",
   954 => x"0000",
   955 => x"0000",
   956 => x"0000",
   957 => x"0000",
   958 => x"0000",
   959 => x"0000",
   960 => x"0000",
   961 => x"0000",
   962 => x"0000",
   963 => x"0000",
   964 => x"0000",
   965 => x"0000",
   966 => x"0000",
   967 => x"0000",
   968 => x"0000",
   969 => x"0000",
   970 => x"0000",
   971 => x"0000",
   972 => x"0000",
   973 => x"0000",
   974 => x"0000",
   975 => x"0000",
   976 => x"0000",
   977 => x"0000",
   978 => x"0000",
   979 => x"0000",
   980 => x"0000",
   981 => x"0000",
   982 => x"0000",
   983 => x"0000",
   984 => x"0000",
   985 => x"0000",
   986 => x"0000",
   987 => x"0000",
   988 => x"0000",
   989 => x"0000",
   990 => x"0000",
   991 => x"0000",
   992 => x"0000",
   993 => x"0000",
   994 => x"0000",
   995 => x"0000",
   996 => x"0000",
   997 => x"0000",
   998 => x"0000",
   999 => x"0000",
  1000 => x"0000",
  1001 => x"0000",
  1002 => x"0000",
  1003 => x"0000",
  1004 => x"0000",
  1005 => x"0000",
  1006 => x"0000",
  1007 => x"0000",
  1008 => x"0000",
  1009 => x"0000",
  1010 => x"0000",
  1011 => x"0000",
  1012 => x"0000",
  1013 => x"0000",
  1014 => x"0000",
  1015 => x"0000",
  1016 => x"0000",
  1017 => x"0000",
  1018 => x"0000",
  1019 => x"0000",
  1020 => x"0000",
  1021 => x"0000",
  1022 => x"0000",
  1023 => x"0000",
  1024 => x"0000",
  1025 => x"0000",
  1026 => x"0000",
  1027 => x"0000",
  1028 => x"0000",
  1029 => x"0000",
  1030 => x"0000",
  1031 => x"0000",
  1032 => x"0000",
  1033 => x"0000",
  1034 => x"0000",
  1035 => x"0000",
  1036 => x"0000",
  1037 => x"0000",
  1038 => x"0000",
  1039 => x"0000",
  1040 => x"0000",
  1041 => x"0000",
  1042 => x"0000",
  1043 => x"0000",
  1044 => x"0000",
  1045 => x"0000",
  1046 => x"0000",
  1047 => x"0000",
  1048 => x"0000",
  1049 => x"0000",
  1050 => x"0000",
  1051 => x"0000",
  1052 => x"0000",
  1053 => x"0000",
  1054 => x"0000",
  1055 => x"0000",
  1056 => x"0000",
  1057 => x"0000",
  1058 => x"0000",
  1059 => x"0000",
  1060 => x"0000",
  1061 => x"0000",
  1062 => x"0000",
  1063 => x"0000",
  1064 => x"0000",
  1065 => x"0000",
  1066 => x"0000",
  1067 => x"0000",
  1068 => x"0000",
  1069 => x"0000",
  1070 => x"0000",
  1071 => x"0000",
  1072 => x"0000",
  1073 => x"0000",
  1074 => x"0000",
  1075 => x"0000",
  1076 => x"0000",
  1077 => x"0000",
  1078 => x"0000",
  1079 => x"0000",
  1080 => x"0000",
  1081 => x"0000",
  1082 => x"0000",
  1083 => x"0000",
  1084 => x"0000",
  1085 => x"0000",
  1086 => x"0000",
  1087 => x"0000",
  1088 => x"0000",
  1089 => x"0000",
  1090 => x"0000",
  1091 => x"0000",
  1092 => x"0000",
  1093 => x"0000",
  1094 => x"0000",
  1095 => x"0000",
  1096 => x"0000",
  1097 => x"0000",
  1098 => x"0000",
  1099 => x"0000",
  1100 => x"0000",
  1101 => x"0000",
  1102 => x"0000",
  1103 => x"0000",
  1104 => x"0000",
  1105 => x"0000",
  1106 => x"0000",
  1107 => x"0000",
  1108 => x"0000",
  1109 => x"0000",
  1110 => x"0000",
  1111 => x"0000",
  1112 => x"0000",
  1113 => x"0000",
  1114 => x"0000",
  1115 => x"0000",
  1116 => x"0000",
  1117 => x"0000",
  1118 => x"0000",
  1119 => x"0000",
  1120 => x"0000",
  1121 => x"0000",
  1122 => x"0000",
  1123 => x"0000",
  1124 => x"0000",
  1125 => x"0000",
  1126 => x"0000",
  1127 => x"0000",
  1128 => x"0000",
  1129 => x"0000",
  1130 => x"0000",
  1131 => x"0000",
  1132 => x"0000",
  1133 => x"0000",
  1134 => x"0000",
  1135 => x"0000",
  1136 => x"0000",
  1137 => x"0000",
  1138 => x"0000",
  1139 => x"0000",
  1140 => x"0000",
  1141 => x"0000",
  1142 => x"0000",
  1143 => x"0000",
  1144 => x"0000",
  1145 => x"0000",
  1146 => x"0000",
  1147 => x"0000",
  1148 => x"0000",
  1149 => x"0000",
  1150 => x"0000",
  1151 => x"0000",
  1152 => x"0000",
  1153 => x"0000",
  1154 => x"0000",
  1155 => x"0000",
  1156 => x"0000",
  1157 => x"0000",
  1158 => x"0000",
  1159 => x"0000",
  1160 => x"0000",
  1161 => x"0000",
  1162 => x"0000",
  1163 => x"0000",
  1164 => x"0000",
  1165 => x"0000",
  1166 => x"0000",
  1167 => x"0000",
  1168 => x"0000",
  1169 => x"0000",
  1170 => x"0000",
  1171 => x"0000",
  1172 => x"0000",
  1173 => x"0000",
  1174 => x"0000",
  1175 => x"0000",
  1176 => x"0000",
  1177 => x"0000",
  1178 => x"0000",
  1179 => x"0000",
  1180 => x"0000",
  1181 => x"0000",
  1182 => x"0000",
  1183 => x"0000",
  1184 => x"0000",
  1185 => x"0000",
  1186 => x"0000",
  1187 => x"0000",
  1188 => x"0000",
  1189 => x"0000",
  1190 => x"0000",
  1191 => x"0000",
  1192 => x"0000",
  1193 => x"0000",
  1194 => x"0000",
  1195 => x"0000",
  1196 => x"0000",
  1197 => x"0000",
  1198 => x"0000",
  1199 => x"0000",
  1200 => x"0000",
  1201 => x"0000",
  1202 => x"0000",
  1203 => x"0000",
  1204 => x"0000",
  1205 => x"0000",
  1206 => x"0000",
  1207 => x"0000",
  1208 => x"0000",
  1209 => x"0000",
  1210 => x"0000",
  1211 => x"0000",
  1212 => x"0000",
  1213 => x"0000",
  1214 => x"0000",
  1215 => x"0000",
  1216 => x"0000",
  1217 => x"0000",
  1218 => x"0000",
  1219 => x"0000",
  1220 => x"0000",
  1221 => x"0000",
  1222 => x"0000",
  1223 => x"0000",
  1224 => x"0000",
  1225 => x"0000",
  1226 => x"0000",
  1227 => x"0000",
  1228 => x"0000",
  1229 => x"0000",
  1230 => x"0000",
  1231 => x"0000",
  1232 => x"0000",
  1233 => x"0000",
  1234 => x"0000",
  1235 => x"0000",
  1236 => x"0000",
  1237 => x"0000",
  1238 => x"0000",
  1239 => x"0000",
  1240 => x"0000",
  1241 => x"0000",
  1242 => x"0000",
  1243 => x"0000",
  1244 => x"0000",
  1245 => x"0000",
  1246 => x"0000",
  1247 => x"0000",
  1248 => x"0000",
  1249 => x"0000",
  1250 => x"0000",
  1251 => x"0000",
  1252 => x"0000",
  1253 => x"0000",
  1254 => x"0000",
  1255 => x"0000",
  1256 => x"0000",
  1257 => x"0000",
  1258 => x"0000",
  1259 => x"0000",
  1260 => x"0000",
  1261 => x"0000",
  1262 => x"0000",
  1263 => x"0000",
  1264 => x"0000",
  1265 => x"0000",
  1266 => x"0000",
  1267 => x"0000",
  1268 => x"0000",
  1269 => x"0000",
  1270 => x"0000",
  1271 => x"0000",
  1272 => x"0000",
  1273 => x"0000",
  1274 => x"0000",
  1275 => x"0000",
  1276 => x"0000",
  1277 => x"0000",
  1278 => x"0000",
  1279 => x"0000",
  1280 => x"0000",
  1281 => x"0000",
  1282 => x"0000",
  1283 => x"0000",
  1284 => x"0000",
  1285 => x"0000",
  1286 => x"0000",
  1287 => x"0000",
  1288 => x"0000",
  1289 => x"0000",
  1290 => x"0000",
  1291 => x"0000",
  1292 => x"0000",
  1293 => x"0000",
  1294 => x"0000",
  1295 => x"0000",
  1296 => x"0000",
  1297 => x"0000",
  1298 => x"0000",
  1299 => x"0000",
  1300 => x"0000",
  1301 => x"0000",
  1302 => x"0000",
  1303 => x"0000",
  1304 => x"0000",
  1305 => x"0000",
  1306 => x"0000",
  1307 => x"0000",
  1308 => x"0000",
  1309 => x"0000",
  1310 => x"0000",
  1311 => x"0000",
  1312 => x"0000",
  1313 => x"0000",
  1314 => x"0000",
  1315 => x"0000",
  1316 => x"0000",
  1317 => x"0000",
  1318 => x"0000",
  1319 => x"0000",
  1320 => x"0000",
  1321 => x"0000",
  1322 => x"0000",
  1323 => x"0000",
  1324 => x"0000",
  1325 => x"0000",
  1326 => x"0000",
  1327 => x"0000",
  1328 => x"0000",
  1329 => x"0000",
  1330 => x"0000",
  1331 => x"0000",
  1332 => x"0000",
  1333 => x"0000",
  1334 => x"0000",
  1335 => x"0000",
  1336 => x"0000",
  1337 => x"0000",
  1338 => x"0000",
  1339 => x"0000",
  1340 => x"0000",
  1341 => x"0000",
  1342 => x"0000",
  1343 => x"0000",
  1344 => x"0000",
  1345 => x"0000",
  1346 => x"0000",
  1347 => x"0000",
  1348 => x"0000",
  1349 => x"0000",
  1350 => x"0000",
  1351 => x"0000",
  1352 => x"0000",
  1353 => x"0000",
  1354 => x"0000",
  1355 => x"0000",
  1356 => x"0000",
  1357 => x"0000",
  1358 => x"0000",
  1359 => x"0000",
  1360 => x"0000",
  1361 => x"0000",
  1362 => x"0000",
  1363 => x"0000",
  1364 => x"0000",
  1365 => x"0000",
  1366 => x"0000",
  1367 => x"0000",
  1368 => x"0000",
  1369 => x"0000",
  1370 => x"0000",
  1371 => x"0000",
  1372 => x"0000",
  1373 => x"0000",
  1374 => x"0000",
  1375 => x"0000",
  1376 => x"0000",
  1377 => x"0000",
  1378 => x"0000",
  1379 => x"0000",
  1380 => x"0000",
  1381 => x"0000",
  1382 => x"0000",
  1383 => x"0000",
  1384 => x"0000",
  1385 => x"0000",
  1386 => x"0000",
  1387 => x"0000",
  1388 => x"0000",
  1389 => x"0000",
  1390 => x"0000",
  1391 => x"0000",
  1392 => x"0000",
  1393 => x"0000",
  1394 => x"0000",
  1395 => x"0000",
  1396 => x"0000",
  1397 => x"0000",
  1398 => x"0000",
  1399 => x"0000",
  1400 => x"0000",
  1401 => x"0000",
  1402 => x"0000",
  1403 => x"0000",
  1404 => x"0000",
  1405 => x"0000",
  1406 => x"0000",
  1407 => x"0000",
  1408 => x"0000",
  1409 => x"0000",
  1410 => x"0000",
  1411 => x"0000",
  1412 => x"0000",
  1413 => x"0000",
  1414 => x"0000",
  1415 => x"0000",
  1416 => x"0000",
  1417 => x"0000",
  1418 => x"0000",
  1419 => x"0000",
  1420 => x"0000",
  1421 => x"0000",
  1422 => x"0000",
  1423 => x"0000",
  1424 => x"0000",
  1425 => x"0000",
  1426 => x"0000",
  1427 => x"0000",
  1428 => x"0000",
  1429 => x"0000",
  1430 => x"0000",
  1431 => x"0000",
  1432 => x"0000",
  1433 => x"0000",
  1434 => x"0000",
  1435 => x"0000",
  1436 => x"0000",
  1437 => x"0000",
  1438 => x"0000",
  1439 => x"0000",
  1440 => x"0000",
  1441 => x"0000",
  1442 => x"0000",
  1443 => x"0000",
  1444 => x"0000",
  1445 => x"0000",
  1446 => x"0000",
  1447 => x"0000",
  1448 => x"0000",
  1449 => x"0000",
  1450 => x"0000",
  1451 => x"0000",
  1452 => x"0000",
  1453 => x"0000",
  1454 => x"0000",
  1455 => x"0000",
  1456 => x"0000",
  1457 => x"0000",
  1458 => x"0000",
  1459 => x"0000",
  1460 => x"0000",
  1461 => x"0000",
  1462 => x"0000",
  1463 => x"0000",
  1464 => x"0000",
  1465 => x"0000",
  1466 => x"0000",
  1467 => x"0000",
  1468 => x"0000",
  1469 => x"0000",
  1470 => x"0000",
  1471 => x"0000",
  1472 => x"0000",
  1473 => x"0000",
  1474 => x"0000",
  1475 => x"0000",
  1476 => x"0000",
  1477 => x"0000",
  1478 => x"0000",
  1479 => x"0000",
  1480 => x"0000",
  1481 => x"0000",
  1482 => x"0000",
  1483 => x"0000",
  1484 => x"0000",
  1485 => x"0000",
  1486 => x"0000",
  1487 => x"0000",
  1488 => x"0000",
  1489 => x"0000",
  1490 => x"0000",
  1491 => x"0000",
  1492 => x"0000",
  1493 => x"0000",
  1494 => x"0000",
  1495 => x"0000",
  1496 => x"0000",
  1497 => x"0000",
  1498 => x"0000",
  1499 => x"0000",
  1500 => x"0000",
  1501 => x"0000",
  1502 => x"0000",
  1503 => x"0000",
  1504 => x"0000",
  1505 => x"0000",
  1506 => x"0000",
  1507 => x"0000",
  1508 => x"0000",
  1509 => x"0000",
  1510 => x"0000",
  1511 => x"0000",
  1512 => x"0000",
  1513 => x"0000",
  1514 => x"0000",
  1515 => x"0000",
  1516 => x"0000",
  1517 => x"0000",
  1518 => x"0000",
  1519 => x"0000",
  1520 => x"0000",
  1521 => x"0000",
  1522 => x"0000",
  1523 => x"0000",
  1524 => x"0000",
  1525 => x"0000",
  1526 => x"0000",
  1527 => x"0000",
  1528 => x"0000",
  1529 => x"0000",
  1530 => x"0000",
  1531 => x"0000",
  1532 => x"0000",
  1533 => x"0000",
  1534 => x"0000",
  1535 => x"0000",
  1536 => x"0000",
  1537 => x"0000",
  1538 => x"0000",
  1539 => x"0000",
  1540 => x"0000",
  1541 => x"0000",
  1542 => x"0000",
  1543 => x"0000",
  1544 => x"0000",
  1545 => x"0000",
  1546 => x"0000",
  1547 => x"0000",
  1548 => x"0000",
  1549 => x"0000",
  1550 => x"0000",
  1551 => x"0000",
  1552 => x"0000",
  1553 => x"0000",
  1554 => x"0000",
  1555 => x"0000",
  1556 => x"0000",
  1557 => x"0000",
  1558 => x"0000",
  1559 => x"0000",
  1560 => x"0000",
  1561 => x"0000",
  1562 => x"0000",
  1563 => x"0000",
  1564 => x"0000",
  1565 => x"0000",
  1566 => x"0000",
  1567 => x"0000",
  1568 => x"0000",
  1569 => x"0000",
  1570 => x"0000",
  1571 => x"0000",
  1572 => x"0000",
  1573 => x"0000",
  1574 => x"0000",
  1575 => x"0000",
  1576 => x"0000",
  1577 => x"0000",
  1578 => x"0000",
  1579 => x"0000",
  1580 => x"0000",
  1581 => x"0000",
  1582 => x"0000",
  1583 => x"0000",
  1584 => x"0000",
  1585 => x"0000",
  1586 => x"0000",
  1587 => x"0000",
  1588 => x"0000",
  1589 => x"0000",
  1590 => x"0000",
  1591 => x"0000",
  1592 => x"0000",
  1593 => x"0000",
  1594 => x"0000",
  1595 => x"0000",
  1596 => x"0000",
  1597 => x"0000",
  1598 => x"0000",
  1599 => x"0000",
  1600 => x"0000",
  1601 => x"0000",
  1602 => x"0000",
  1603 => x"0000",
  1604 => x"0000",
  1605 => x"0000",
  1606 => x"0000",
  1607 => x"0000",
  1608 => x"0000",
  1609 => x"0000",
  1610 => x"0000",
  1611 => x"0000",
  1612 => x"0000",
  1613 => x"0000",
  1614 => x"0000",
  1615 => x"0000",
  1616 => x"0000",
  1617 => x"0000",
  1618 => x"0000",
  1619 => x"0000",
  1620 => x"0000",
  1621 => x"0000",
  1622 => x"0000",
  1623 => x"0000",
  1624 => x"0000",
  1625 => x"0000",
  1626 => x"0000",
  1627 => x"0000",
  1628 => x"0000",
  1629 => x"0000",
  1630 => x"0000",
  1631 => x"0000",
  1632 => x"0000",
  1633 => x"0000",
  1634 => x"0000",
  1635 => x"0000",
  1636 => x"0000",
  1637 => x"0000",
  1638 => x"0000",
  1639 => x"0000",
  1640 => x"0000",
  1641 => x"0000",
  1642 => x"0000",
  1643 => x"0000",
  1644 => x"0000",
  1645 => x"0000",
  1646 => x"0000",
  1647 => x"0000",
  1648 => x"0000",
  1649 => x"0000",
  1650 => x"0000",
  1651 => x"0000",
  1652 => x"0000",
  1653 => x"0000",
  1654 => x"0000",
  1655 => x"0000",
  1656 => x"0000",
  1657 => x"0000",
  1658 => x"0000",
  1659 => x"0000",
  1660 => x"0000",
  1661 => x"0000",
  1662 => x"0000",
  1663 => x"0000",
  1664 => x"0000",
  1665 => x"0000",
  1666 => x"0000",
  1667 => x"0000",
  1668 => x"0000",
  1669 => x"0000",
  1670 => x"0000",
  1671 => x"0000",
  1672 => x"0000",
  1673 => x"0000",
  1674 => x"0000",
  1675 => x"0000",
  1676 => x"0000",
  1677 => x"0000",
  1678 => x"0000",
  1679 => x"0000",
  1680 => x"0000",
  1681 => x"0000",
  1682 => x"0000",
  1683 => x"0000",
  1684 => x"0000",
  1685 => x"0000",
  1686 => x"0000",
  1687 => x"0000",
  1688 => x"0000",
  1689 => x"0000",
  1690 => x"0000",
  1691 => x"0000",
  1692 => x"0000",
  1693 => x"0000",
  1694 => x"0000",
  1695 => x"0000",
  1696 => x"0000",
  1697 => x"0000",
  1698 => x"0000",
  1699 => x"0000",
  1700 => x"0000",
  1701 => x"0000",
  1702 => x"0000",
  1703 => x"0000",
  1704 => x"0000",
  1705 => x"0000",
  1706 => x"0000",
  1707 => x"0000",
  1708 => x"0000",
  1709 => x"0000",
  1710 => x"0000",
  1711 => x"0000",
  1712 => x"0000",
  1713 => x"0000",
  1714 => x"0000",
  1715 => x"0000",
  1716 => x"0000",
  1717 => x"0000",
  1718 => x"0000",
  1719 => x"0000",
  1720 => x"0000",
  1721 => x"0000",
  1722 => x"0000",
  1723 => x"0000",
  1724 => x"0000",
  1725 => x"0000",
  1726 => x"0000",
  1727 => x"0000",
  1728 => x"0000",
  1729 => x"0000",
  1730 => x"0000",
  1731 => x"0000",
  1732 => x"0000",
  1733 => x"0000",
  1734 => x"0000",
  1735 => x"0000",
  1736 => x"0000",
  1737 => x"0000",
  1738 => x"0000",
  1739 => x"0000",
  1740 => x"0000",
  1741 => x"0000",
  1742 => x"0000",
  1743 => x"0000",
  1744 => x"0000",
  1745 => x"0000",
  1746 => x"0000",
  1747 => x"0000",
  1748 => x"0000",
  1749 => x"0000",
  1750 => x"0000",
  1751 => x"0000",
  1752 => x"0000",
  1753 => x"0000",
  1754 => x"0000",
  1755 => x"0000",
  1756 => x"0000",
  1757 => x"0000",
  1758 => x"0000",
  1759 => x"0000",
  1760 => x"0000",
  1761 => x"0000",
  1762 => x"0000",
  1763 => x"0000",
  1764 => x"0000",
  1765 => x"0000",
  1766 => x"0000",
  1767 => x"0000",
  1768 => x"0000",
  1769 => x"0000",
  1770 => x"0000",
  1771 => x"0000",
  1772 => x"0000",
  1773 => x"0000",
  1774 => x"0000",
  1775 => x"0000",
  1776 => x"0000",
  1777 => x"0000",
  1778 => x"0000",
  1779 => x"0000",
  1780 => x"0000",
  1781 => x"0000",
  1782 => x"0000",
  1783 => x"0000",
  1784 => x"0000",
  1785 => x"0000",
  1786 => x"0000",
  1787 => x"0000",
  1788 => x"0000",
  1789 => x"0000",
  1790 => x"0000",
  1791 => x"0000",
  1792 => x"0000",
  1793 => x"0000",
  1794 => x"0000",
  1795 => x"0000",
  1796 => x"0000",
  1797 => x"0000",
  1798 => x"0000",
  1799 => x"0000",
  1800 => x"0000",
  1801 => x"0000",
  1802 => x"0000",
  1803 => x"0000",
  1804 => x"0000",
  1805 => x"0000",
  1806 => x"0000",
  1807 => x"0000",
  1808 => x"0000",
  1809 => x"0000",
  1810 => x"0000",
  1811 => x"0000",
  1812 => x"0000",
  1813 => x"0000",
  1814 => x"0000",
  1815 => x"0000",
  1816 => x"0000",
  1817 => x"0000",
  1818 => x"0000",
  1819 => x"0000",
  1820 => x"0000",
  1821 => x"0000",
  1822 => x"0000",
  1823 => x"0000",
  1824 => x"0000",
  1825 => x"0000",
  1826 => x"0000",
  1827 => x"0000",
  1828 => x"0000",
  1829 => x"0000",
  1830 => x"0000",
  1831 => x"0000",
  1832 => x"0000",
  1833 => x"0000",
  1834 => x"0000",
  1835 => x"0000",
  1836 => x"0000",
  1837 => x"0000",
  1838 => x"0000",
  1839 => x"0000",
  1840 => x"0000",
  1841 => x"0000",
  1842 => x"0000",
  1843 => x"0000",
  1844 => x"0000",
  1845 => x"0000",
  1846 => x"0000",
  1847 => x"0000",
  1848 => x"0000",
  1849 => x"0000",
  1850 => x"0000",
  1851 => x"0000",
  1852 => x"0000",
  1853 => x"0000",
  1854 => x"0000",
  1855 => x"0000",
  1856 => x"0000",
  1857 => x"0000",
  1858 => x"0000",
  1859 => x"0000",
  1860 => x"0000",
  1861 => x"0000",
  1862 => x"0000",
  1863 => x"0000",
  1864 => x"0000",
  1865 => x"0000",
  1866 => x"0000",
  1867 => x"0000",
  1868 => x"0000",
  1869 => x"0000",
  1870 => x"0000",
  1871 => x"0000",
  1872 => x"0000",
  1873 => x"0000",
  1874 => x"0000",
  1875 => x"0000",
  1876 => x"0000",
  1877 => x"0000",
  1878 => x"0000",
  1879 => x"0000",
  1880 => x"0000",
  1881 => x"0000",
  1882 => x"0000",
  1883 => x"0000",
  1884 => x"0000",
  1885 => x"0000",
  1886 => x"0000",
  1887 => x"0000",
  1888 => x"0000",
  1889 => x"0000",
  1890 => x"0000",
  1891 => x"0000",
  1892 => x"0000",
  1893 => x"0000",
  1894 => x"0000",
  1895 => x"0000",
  1896 => x"0000",
  1897 => x"0000",
  1898 => x"0000",
  1899 => x"0000",
  1900 => x"0000",
  1901 => x"0000",
  1902 => x"0000",
  1903 => x"0000",
  1904 => x"0000",
  1905 => x"0000",
  1906 => x"0000",
  1907 => x"0000",
  1908 => x"0000",
  1909 => x"0000",
  1910 => x"0000",
  1911 => x"0000",
  1912 => x"0000",
  1913 => x"0000",
  1914 => x"0000",
  1915 => x"0000",
  1916 => x"0000",
  1917 => x"0000",
  1918 => x"0000",
  1919 => x"0000",
  1920 => x"0000",
  1921 => x"0000",
  1922 => x"0000",
  1923 => x"0000",
  1924 => x"0000",
  1925 => x"0000",
  1926 => x"0000",
  1927 => x"0000",
  1928 => x"0000",
  1929 => x"0000",
  1930 => x"0000",
  1931 => x"0000",
  1932 => x"0000",
  1933 => x"0000",
  1934 => x"0000",
  1935 => x"0000",
  1936 => x"0000",
  1937 => x"0000",
  1938 => x"0000",
  1939 => x"0000",
  1940 => x"0000",
  1941 => x"0000",
  1942 => x"0000",
  1943 => x"0000",
  1944 => x"0000",
  1945 => x"0000",
  1946 => x"0000",
  1947 => x"0000",
  1948 => x"0000",
  1949 => x"0000",
  1950 => x"0000",
  1951 => x"0000",
  1952 => x"0000",
  1953 => x"0000",
  1954 => x"0000",
  1955 => x"0000",
  1956 => x"0000",
  1957 => x"0000",
  1958 => x"0000",
  1959 => x"0000",
  1960 => x"0000",
  1961 => x"0000",
  1962 => x"0000",
  1963 => x"0000",
  1964 => x"0000",
  1965 => x"0000",
  1966 => x"0000",
  1967 => x"0000",
  1968 => x"0000",
  1969 => x"0000",
  1970 => x"0000",
  1971 => x"0000",
  1972 => x"0000",
  1973 => x"0000",
  1974 => x"0000",
  1975 => x"0000",
  1976 => x"0000",
  1977 => x"0000",
  1978 => x"0000",
  1979 => x"0000",
  1980 => x"0000",
  1981 => x"0000",
  1982 => x"0000",
  1983 => x"0000",
  1984 => x"0000",
  1985 => x"0000",
  1986 => x"0000",
  1987 => x"0000",
  1988 => x"0000",
  1989 => x"0000",
  1990 => x"0000",
  1991 => x"0000",
  1992 => x"0000",
  1993 => x"0000",
  1994 => x"0000",
  1995 => x"0000",
  1996 => x"0000",
  1997 => x"0000",
  1998 => x"0000",
  1999 => x"0000",
  2000 => x"0000",
  2001 => x"0000",
  2002 => x"0000",
  2003 => x"0000",
  2004 => x"0000",
  2005 => x"0000",
  2006 => x"0000",
  2007 => x"0000",
  2008 => x"0000",
  2009 => x"0000",
  2010 => x"0000",
  2011 => x"0000",
  2012 => x"0000",
  2013 => x"0000",
  2014 => x"0000",
  2015 => x"0000",
  2016 => x"0000",
  2017 => x"0000",
  2018 => x"0000",
  2019 => x"0000",
  2020 => x"0000",
  2021 => x"0000",
  2022 => x"0000",
  2023 => x"0000",
  2024 => x"0000",
  2025 => x"0000",
  2026 => x"0000",
  2027 => x"0000",
  2028 => x"0000",
  2029 => x"0000",
  2030 => x"0000",
  2031 => x"0000",
  2032 => x"0000",
  2033 => x"0000",
  2034 => x"0000",
  2035 => x"0000",
  2036 => x"0000",
  2037 => x"0000",
  2038 => x"0000",
  2039 => x"0000",
  2040 => x"0000",
  2041 => x"0000",
  2042 => x"0000",
  2043 => x"0000",
  2044 => x"0000",
  2045 => x"0000",
  2046 => x"0000",
  2047 => x"0000",
  2048 => x"0000",
  2049 => x"0000",
  2050 => x"0000",
  2051 => x"0000",
  2052 => x"0000",
  2053 => x"0000",
  2054 => x"0000",
  2055 => x"0000",
  2056 => x"0000",
  2057 => x"0000",
  2058 => x"0000",
  2059 => x"0000",
  2060 => x"0000",
  2061 => x"0000",
  2062 => x"0000",
  2063 => x"0000",
  2064 => x"0000",
  2065 => x"0000",
  2066 => x"0000",
  2067 => x"0000",
  2068 => x"0000",
  2069 => x"0000",
  2070 => x"0000",
  2071 => x"0000",
  2072 => x"0000",
  2073 => x"0000",
  2074 => x"0000",
  2075 => x"0000",
  2076 => x"0000",
  2077 => x"0000",
  2078 => x"0000",
  2079 => x"0000",
  2080 => x"0000",
  2081 => x"0000",
  2082 => x"0000",
  2083 => x"0000",
  2084 => x"0000",
  2085 => x"0000",
  2086 => x"0000",
  2087 => x"0000",
  2088 => x"0000",
  2089 => x"0000",
  2090 => x"0000",
  2091 => x"0000",
  2092 => x"0000",
  2093 => x"0000",
  2094 => x"0000",
  2095 => x"0000",
  2096 => x"0000",
  2097 => x"0000",
  2098 => x"0000",
  2099 => x"0000",
  2100 => x"0000",
  2101 => x"0000",
  2102 => x"0000",
  2103 => x"0000",
  2104 => x"0000",
  2105 => x"0000",
  2106 => x"0000",
  2107 => x"0000",
  2108 => x"0000",
  2109 => x"0000",
  2110 => x"0000",
  2111 => x"0000",
  2112 => x"0000",
  2113 => x"0000",
  2114 => x"0000",
  2115 => x"0000",
  2116 => x"0000",
  2117 => x"0000",
  2118 => x"0000",
  2119 => x"0000",
  2120 => x"0000",
  2121 => x"0000",
  2122 => x"0000",
  2123 => x"0000",
  2124 => x"0000",
  2125 => x"0000",
  2126 => x"0000",
  2127 => x"0000",
  2128 => x"0000",
  2129 => x"0000",
  2130 => x"0000",
  2131 => x"0000",
  2132 => x"0000",
  2133 => x"0000",
  2134 => x"0000",
  2135 => x"0000",
  2136 => x"0000",
  2137 => x"0000",
  2138 => x"0000",
  2139 => x"0000",
  2140 => x"0000",
  2141 => x"0000",
  2142 => x"0000",
  2143 => x"0000",
  2144 => x"0000",
  2145 => x"0000",
  2146 => x"0000",
  2147 => x"0000",
  2148 => x"0000",
  2149 => x"0000",
  2150 => x"0000",
  2151 => x"0000",
  2152 => x"0000",
  2153 => x"0000",
  2154 => x"0000",
  2155 => x"0000",
  2156 => x"0000",
  2157 => x"0000",
  2158 => x"0000",
  2159 => x"0000",
  2160 => x"0000",
  2161 => x"0000",
  2162 => x"0000",
  2163 => x"0000",
  2164 => x"0000",
  2165 => x"0000",
  2166 => x"0000",
  2167 => x"0000",
  2168 => x"0000",
  2169 => x"0000",
  2170 => x"0000",
  2171 => x"0000",
  2172 => x"0000",
  2173 => x"0000",
  2174 => x"0000",
  2175 => x"0000",
  2176 => x"0000",
  2177 => x"0000",
  2178 => x"0000",
  2179 => x"0000",
  2180 => x"0000",
  2181 => x"0000",
  2182 => x"0000",
  2183 => x"0000",
  2184 => x"0000",
  2185 => x"0000",
  2186 => x"0000",
  2187 => x"0000",
  2188 => x"0000",
  2189 => x"0000",
  2190 => x"0000",
  2191 => x"0000",
  2192 => x"0000",
  2193 => x"0000",
  2194 => x"0000",
  2195 => x"0000",
  2196 => x"0000",
  2197 => x"0000",
  2198 => x"0000",
  2199 => x"0000",
  2200 => x"0000",
  2201 => x"0000",
  2202 => x"0000",
  2203 => x"0000",
  2204 => x"0000",
  2205 => x"0000",
  2206 => x"0000",
  2207 => x"0000",
  2208 => x"0000",
  2209 => x"0000",
  2210 => x"0000",
  2211 => x"0000",
  2212 => x"0000",
  2213 => x"0000",
  2214 => x"0000",
  2215 => x"0000",
  2216 => x"0000",
  2217 => x"0000",
  2218 => x"0000",
  2219 => x"0000",
  2220 => x"0000",
  2221 => x"0000",
  2222 => x"0000",
  2223 => x"0000",
  2224 => x"0000",
  2225 => x"0000",
  2226 => x"0000",
  2227 => x"0000",
  2228 => x"0000",
  2229 => x"0000",
  2230 => x"0000",
  2231 => x"0000",
  2232 => x"0000",
  2233 => x"0000",
  2234 => x"0000",
  2235 => x"0000",
  2236 => x"0000",
  2237 => x"0000",
  2238 => x"0000",
  2239 => x"0000",
  2240 => x"0000",
  2241 => x"0000",
  2242 => x"0000",
  2243 => x"0000",
  2244 => x"0000",
  2245 => x"0000",
  2246 => x"0000",
  2247 => x"0000",
  2248 => x"0000",
  2249 => x"0000",
  2250 => x"0000",
  2251 => x"0000",
  2252 => x"0000",
  2253 => x"0000",
  2254 => x"0000",
  2255 => x"0000",
  2256 => x"0000",
  2257 => x"0000",
  2258 => x"0000",
  2259 => x"0000",
  2260 => x"0000",
  2261 => x"0000",
  2262 => x"0000",
  2263 => x"0000",
  2264 => x"0000",
  2265 => x"0000",
  2266 => x"0000",
  2267 => x"0000",
  2268 => x"0000",
  2269 => x"0000",
  2270 => x"0000",
  2271 => x"0000",
  2272 => x"0000",
  2273 => x"0000",
  2274 => x"0000",
  2275 => x"0000",
  2276 => x"0000",
  2277 => x"0000",
  2278 => x"0000",
  2279 => x"0000",
  2280 => x"0000",
  2281 => x"0000",
  2282 => x"0000",
  2283 => x"0000",
  2284 => x"0000",
  2285 => x"0000",
  2286 => x"0000",
  2287 => x"0000",
  2288 => x"0000",
  2289 => x"0000",
  2290 => x"0000",
  2291 => x"0000",
  2292 => x"0000",
  2293 => x"0000",
  2294 => x"0000",
  2295 => x"0000",
  2296 => x"0000",
  2297 => x"0000",
  2298 => x"0000",
  2299 => x"0000",
  2300 => x"0000",
  2301 => x"0000",
  2302 => x"0000",
  2303 => x"0000",
  2304 => x"0000",
  2305 => x"0000",
  2306 => x"0000",
  2307 => x"0000",
  2308 => x"0000",
  2309 => x"0000",
  2310 => x"0000",
  2311 => x"0000",
  2312 => x"0000",
  2313 => x"0000",
  2314 => x"0000",
  2315 => x"0000",
  2316 => x"0000",
  2317 => x"0000",
  2318 => x"0000",
  2319 => x"0000",
  2320 => x"0000",
  2321 => x"0000",
  2322 => x"0000",
  2323 => x"0000",
  2324 => x"0000",
  2325 => x"0000",
  2326 => x"0000",
  2327 => x"0000",
  2328 => x"0000",
  2329 => x"0000",
  2330 => x"0000",
  2331 => x"0000",
  2332 => x"0000",
  2333 => x"0000",
  2334 => x"0000",
  2335 => x"0000",
  2336 => x"0000",
  2337 => x"0000",
  2338 => x"0000",
  2339 => x"0000",
  2340 => x"0000",
  2341 => x"0000",
  2342 => x"0000",
  2343 => x"0000",
  2344 => x"0000",
  2345 => x"0000",
  2346 => x"0000",
  2347 => x"0000",
  2348 => x"0000",
  2349 => x"0000",
  2350 => x"0000",
  2351 => x"0000",
  2352 => x"0000",
  2353 => x"0000",
  2354 => x"0000",
  2355 => x"0000",
  2356 => x"0000",
  2357 => x"0000",
  2358 => x"0000",
  2359 => x"0000",
  2360 => x"0000",
  2361 => x"0000",
  2362 => x"0000",
  2363 => x"0000",
  2364 => x"0000",
  2365 => x"0000",
  2366 => x"0000",
  2367 => x"0000",
  2368 => x"0000",
  2369 => x"0000",
  2370 => x"0000",
  2371 => x"0000",
  2372 => x"0000",
  2373 => x"0000",
  2374 => x"0000",
  2375 => x"0000",
  2376 => x"0000",
  2377 => x"0000",
  2378 => x"0000",
  2379 => x"0000",
  2380 => x"0000",
  2381 => x"0000",
  2382 => x"0000",
  2383 => x"0000",
  2384 => x"0000",
  2385 => x"0000",
  2386 => x"0000",
  2387 => x"0000",
  2388 => x"0000",
  2389 => x"0000",
  2390 => x"0000",
  2391 => x"0000",
  2392 => x"0000",
  2393 => x"0000",
  2394 => x"0000",
  2395 => x"0000",
  2396 => x"0000",
  2397 => x"0000",
  2398 => x"0000",
  2399 => x"0000",
  2400 => x"0000",
  2401 => x"0000",
  2402 => x"0000",
  2403 => x"0000",
  2404 => x"0000",
  2405 => x"0000",
  2406 => x"0000",
  2407 => x"0000",
  2408 => x"0000",
  2409 => x"0000",
  2410 => x"0000",
  2411 => x"0000",
  2412 => x"0000",
  2413 => x"0000",
  2414 => x"0000",
  2415 => x"0000",
  2416 => x"0000",
  2417 => x"0000",
  2418 => x"0000",
  2419 => x"0000",
  2420 => x"0000",
  2421 => x"0000",
  2422 => x"0000",
  2423 => x"0000",
  2424 => x"0000",
  2425 => x"0000",
  2426 => x"0000",
  2427 => x"0000",
  2428 => x"0000",
  2429 => x"0000",
  2430 => x"0000",
  2431 => x"0000",
  2432 => x"0000",
  2433 => x"0000",
  2434 => x"0000",
  2435 => x"0000",
  2436 => x"0000",
  2437 => x"0000",
  2438 => x"0000",
  2439 => x"0000",
  2440 => x"0000",
  2441 => x"0000",
  2442 => x"0000",
  2443 => x"0000",
  2444 => x"0000",
  2445 => x"0000",
  2446 => x"0000",
  2447 => x"0000",
  2448 => x"0000",
  2449 => x"0000",
  2450 => x"0000",
  2451 => x"0000",
  2452 => x"0000",
  2453 => x"0000",
  2454 => x"0000",
  2455 => x"0000",
  2456 => x"0000",
  2457 => x"0000",
  2458 => x"0000",
  2459 => x"0000",
  2460 => x"0000",
  2461 => x"0000",
  2462 => x"0000",
  2463 => x"0000",
  2464 => x"0000",
  2465 => x"0000",
  2466 => x"0000",
  2467 => x"0000",
  2468 => x"0000",
  2469 => x"0000",
  2470 => x"0000",
  2471 => x"0000",
  2472 => x"0000",
  2473 => x"0000",
  2474 => x"0000",
  2475 => x"0000",
  2476 => x"0000",
  2477 => x"0000",
  2478 => x"0000",
  2479 => x"0000",
  2480 => x"0000",
  2481 => x"0000",
  2482 => x"0000",
  2483 => x"0000",
  2484 => x"0000",
  2485 => x"0000",
  2486 => x"0000",
  2487 => x"0000",
  2488 => x"0000",
  2489 => x"0000",
  2490 => x"0000",
  2491 => x"0000",
  2492 => x"0000",
  2493 => x"0000",
  2494 => x"0000",
  2495 => x"0000",
  2496 => x"0000",
  2497 => x"0000",
  2498 => x"0000",
  2499 => x"0000",
  2500 => x"0000",
  2501 => x"0000",
  2502 => x"0000",
  2503 => x"0000",
  2504 => x"0000",
  2505 => x"0000",
  2506 => x"0000",
  2507 => x"0000",
  2508 => x"0000",
  2509 => x"0000",
  2510 => x"0000",
  2511 => x"0000",
  2512 => x"0000",
  2513 => x"0000",
  2514 => x"0000",
  2515 => x"0000",
  2516 => x"0000",
  2517 => x"0000",
  2518 => x"0000",
  2519 => x"0000",
  2520 => x"0000",
  2521 => x"0000",
  2522 => x"0000",
  2523 => x"0000",
  2524 => x"0000",
  2525 => x"0000",
  2526 => x"0000",
  2527 => x"0000",
  2528 => x"0000",
  2529 => x"0000",
  2530 => x"0000",
  2531 => x"0000",
  2532 => x"0000",
  2533 => x"0000",
  2534 => x"0000",
  2535 => x"0000",
  2536 => x"0000",
  2537 => x"0000",
  2538 => x"0000",
  2539 => x"0000",
  2540 => x"0000",
  2541 => x"0000",
  2542 => x"0000",
  2543 => x"0000",
  2544 => x"0000",
  2545 => x"0000",
  2546 => x"0000",
  2547 => x"0000",
  2548 => x"0000",
  2549 => x"0000",
  2550 => x"0000",
  2551 => x"0000",
  2552 => x"0000",
  2553 => x"0000",
  2554 => x"0000",
  2555 => x"0000",
  2556 => x"0000",
  2557 => x"0000",
  2558 => x"0000",
  2559 => x"0000",
  2560 => x"0000",
  2561 => x"0000",
  2562 => x"0000",
  2563 => x"0000",
  2564 => x"0000",
  2565 => x"0000",
  2566 => x"0000",
  2567 => x"0000",
  2568 => x"0000",
  2569 => x"0000",
  2570 => x"0000",
  2571 => x"0000",
  2572 => x"0000",
  2573 => x"0000",
  2574 => x"0000",
  2575 => x"0000",
  2576 => x"0000",
  2577 => x"0000",
  2578 => x"0000",
  2579 => x"0000",
  2580 => x"0000",
  2581 => x"0000",
  2582 => x"0000",
  2583 => x"0000",
  2584 => x"0000",
  2585 => x"0000",
  2586 => x"0000",
  2587 => x"0000",
  2588 => x"0000",
  2589 => x"0000",
  2590 => x"0000",
  2591 => x"0000",
  2592 => x"0000",
  2593 => x"0000",
  2594 => x"0000",
  2595 => x"0000",
  2596 => x"0000",
  2597 => x"0000",
  2598 => x"0000",
  2599 => x"0000",
  2600 => x"0000",
  2601 => x"0000",
  2602 => x"0000",
  2603 => x"0000",
  2604 => x"0000",
  2605 => x"0000",
  2606 => x"0000",
  2607 => x"0000",
  2608 => x"0000",
  2609 => x"0000",
  2610 => x"0000",
  2611 => x"0000",
  2612 => x"0000",
  2613 => x"0000",
  2614 => x"0000",
  2615 => x"0000",
  2616 => x"0000",
  2617 => x"0000",
  2618 => x"0000",
  2619 => x"0000",
  2620 => x"0000",
  2621 => x"0000",
  2622 => x"0000",
  2623 => x"0000",
  2624 => x"0000",
  2625 => x"0000",
  2626 => x"0000",
  2627 => x"0000",
  2628 => x"0000",
  2629 => x"0000",
  2630 => x"0000",
  2631 => x"0000",
  2632 => x"0000",
  2633 => x"0000",
  2634 => x"0000",
  2635 => x"0000",
  2636 => x"0000",
  2637 => x"0000",
  2638 => x"0000",
  2639 => x"0000",
  2640 => x"0000",
  2641 => x"0000",
  2642 => x"0000",
  2643 => x"0000",
  2644 => x"0000",
  2645 => x"0000",
  2646 => x"0000",
  2647 => x"0000",
  2648 => x"0000",
  2649 => x"0000",
  2650 => x"0000",
  2651 => x"0000",
  2652 => x"0000",
  2653 => x"0000",
  2654 => x"0000",
  2655 => x"0000",
  2656 => x"0000",
  2657 => x"0000",
  2658 => x"0000",
  2659 => x"0000",
  2660 => x"0000",
  2661 => x"0000",
  2662 => x"0000",
  2663 => x"0000",
  2664 => x"0000",
  2665 => x"0000",
  2666 => x"0000",
  2667 => x"0000",
  2668 => x"0000",
  2669 => x"0000",
  2670 => x"0000",
  2671 => x"0000",
  2672 => x"0000",
  2673 => x"0000",
  2674 => x"0000",
  2675 => x"0000",
  2676 => x"0000",
  2677 => x"0000",
  2678 => x"0000",
  2679 => x"0000",
  2680 => x"0000",
  2681 => x"0000",
  2682 => x"0000",
  2683 => x"0000",
  2684 => x"0000",
  2685 => x"0000",
  2686 => x"0000",
  2687 => x"0000",
  2688 => x"0000",
  2689 => x"0000",
  2690 => x"0000",
  2691 => x"0000",
  2692 => x"0000",
  2693 => x"0000",
  2694 => x"0000",
  2695 => x"0000",
  2696 => x"0000",
  2697 => x"0000",
  2698 => x"0000",
  2699 => x"0000",
  2700 => x"0000",
  2701 => x"0000",
  2702 => x"0000",
  2703 => x"0000",
  2704 => x"0000",
  2705 => x"0000",
  2706 => x"0000",
  2707 => x"0000",
  2708 => x"0000",
  2709 => x"0000",
  2710 => x"0000",
  2711 => x"0000",
  2712 => x"0000",
  2713 => x"0000",
  2714 => x"0000",
  2715 => x"0000",
  2716 => x"0000",
  2717 => x"0000",
  2718 => x"0000",
  2719 => x"0000",
  2720 => x"0000",
  2721 => x"0000",
  2722 => x"0000",
  2723 => x"0000",
  2724 => x"0000",
  2725 => x"0000",
  2726 => x"0000",
  2727 => x"0000",
  2728 => x"0000",
  2729 => x"0000",
  2730 => x"0000",
  2731 => x"0000",
  2732 => x"0000",
  2733 => x"0000",
  2734 => x"0000",
  2735 => x"0000",
  2736 => x"0000",
  2737 => x"0000",
  2738 => x"0000",
  2739 => x"0000",
  2740 => x"0000",
  2741 => x"0000",
  2742 => x"0000",
  2743 => x"0000",
  2744 => x"0000",
  2745 => x"0000",
  2746 => x"0000",
  2747 => x"0000",
  2748 => x"0000",
  2749 => x"0000",
  2750 => x"0000",
  2751 => x"0000",
  2752 => x"0000",
  2753 => x"0000",
  2754 => x"0000",
  2755 => x"0000",
  2756 => x"0000",
  2757 => x"0000",
  2758 => x"0000",
  2759 => x"0000",
  2760 => x"0000",
  2761 => x"0000",
  2762 => x"0000",
  2763 => x"0000",
  2764 => x"0000",
  2765 => x"0000",
  2766 => x"0000",
  2767 => x"0000",
  2768 => x"0000",
  2769 => x"0000",
  2770 => x"0000",
  2771 => x"0000",
  2772 => x"0000",
  2773 => x"0000",
  2774 => x"0000",
  2775 => x"0000",
  2776 => x"0000",
  2777 => x"0000",
  2778 => x"0000",
  2779 => x"0000",
  2780 => x"0000",
  2781 => x"0000",
  2782 => x"0000",
  2783 => x"0000",
  2784 => x"0000",
  2785 => x"0000",
  2786 => x"0000",
  2787 => x"0000",
  2788 => x"0000",
  2789 => x"0000",
  2790 => x"0000",
  2791 => x"0000",
  2792 => x"0000",
  2793 => x"0000",
  2794 => x"0000",
  2795 => x"0000",
  2796 => x"0000",
  2797 => x"0000",
  2798 => x"0000",
  2799 => x"0000",
  2800 => x"0000",
  2801 => x"0000",
  2802 => x"0000",
  2803 => x"0000",
  2804 => x"0000",
  2805 => x"0000",
  2806 => x"0000",
  2807 => x"0000",
  2808 => x"0000",
  2809 => x"0000",
  2810 => x"0000",
  2811 => x"0000",
  2812 => x"0000",
  2813 => x"0000",
  2814 => x"0000",
  2815 => x"0000",
  2816 => x"0000",
  2817 => x"0000",
  2818 => x"0000",
  2819 => x"0000",
  2820 => x"0000",
  2821 => x"0000",
  2822 => x"0000",
  2823 => x"0000",
  2824 => x"0000",
  2825 => x"0000",
  2826 => x"0000",
  2827 => x"0000",
  2828 => x"0000",
  2829 => x"0000",
  2830 => x"0000",
  2831 => x"0000",
  2832 => x"0000",
  2833 => x"0000",
  2834 => x"0000",
  2835 => x"0000",
  2836 => x"0000",
  2837 => x"0000",
  2838 => x"0000",
  2839 => x"0000",
  2840 => x"0000",
  2841 => x"0000",
  2842 => x"0000",
  2843 => x"0000",
  2844 => x"0000",
  2845 => x"0000",
  2846 => x"0000",
  2847 => x"0000",
  2848 => x"0000",
  2849 => x"0000",
  2850 => x"0000",
  2851 => x"0000",
  2852 => x"0000",
  2853 => x"0000",
  2854 => x"0000",
  2855 => x"0000",
  2856 => x"0000",
  2857 => x"0000",
  2858 => x"0000",
  2859 => x"0000",
  2860 => x"0000",
  2861 => x"0000",
  2862 => x"0000",
  2863 => x"0000",
  2864 => x"0000",
  2865 => x"0000",
  2866 => x"0000",
  2867 => x"0000",
  2868 => x"0000",
  2869 => x"0000",
  2870 => x"0000",
  2871 => x"0000",
  2872 => x"0000",
  2873 => x"0000",
  2874 => x"0000",
  2875 => x"0000",
  2876 => x"0000",
  2877 => x"0000",
  2878 => x"0000",
  2879 => x"0000",
  2880 => x"0000",
  2881 => x"0000",
  2882 => x"0000",
  2883 => x"0000",
  2884 => x"0000",
  2885 => x"0000",
  2886 => x"0000",
  2887 => x"0000",
  2888 => x"0000",
  2889 => x"0000",
  2890 => x"0000",
  2891 => x"0000",
  2892 => x"0000",
  2893 => x"0000",
  2894 => x"0000",
  2895 => x"0000",
  2896 => x"0000",
  2897 => x"0000",
  2898 => x"0000",
  2899 => x"0000",
  2900 => x"0000",
  2901 => x"0000",
  2902 => x"0000",
  2903 => x"0000",
  2904 => x"0000",
  2905 => x"0000",
  2906 => x"0000",
  2907 => x"0000",
  2908 => x"0000",
  2909 => x"0000",
  2910 => x"0000",
  2911 => x"0000",
  2912 => x"0000",
  2913 => x"0000",
  2914 => x"0000",
  2915 => x"0000",
  2916 => x"0000",
  2917 => x"0000",
  2918 => x"0000",
  2919 => x"0000",
  2920 => x"0000",
  2921 => x"0000",
  2922 => x"0000",
  2923 => x"0000",
  2924 => x"0000",
  2925 => x"0000",
  2926 => x"0000",
  2927 => x"0000",
  2928 => x"0000",
  2929 => x"0000",
  2930 => x"0000",
  2931 => x"0000",
  2932 => x"0000",
  2933 => x"0000",
  2934 => x"0000",
  2935 => x"0000",
  2936 => x"0000",
  2937 => x"0000",
  2938 => x"0000",
  2939 => x"0000",
  2940 => x"0000",
  2941 => x"0000",
  2942 => x"0000",
  2943 => x"0000",
  2944 => x"0000",
  2945 => x"0000",
  2946 => x"0000",
  2947 => x"0000",
  2948 => x"0000",
  2949 => x"0000",
  2950 => x"0000",
  2951 => x"0000",
  2952 => x"0000",
  2953 => x"0000",
  2954 => x"0000",
  2955 => x"0000",
  2956 => x"0000",
  2957 => x"0000",
  2958 => x"0000",
  2959 => x"0000",
  2960 => x"0000",
  2961 => x"0000",
  2962 => x"0000",
  2963 => x"0000",
  2964 => x"0000",
  2965 => x"0000",
  2966 => x"0000",
  2967 => x"0000",
  2968 => x"0000",
  2969 => x"0000",
  2970 => x"0000",
  2971 => x"0000",
  2972 => x"0000",
  2973 => x"0000",
  2974 => x"0000",
  2975 => x"0000",
  2976 => x"0000",
  2977 => x"0000",
  2978 => x"0000",
  2979 => x"0000",
  2980 => x"0000",
  2981 => x"0000",
  2982 => x"0000",
  2983 => x"0000",
  2984 => x"0000",
  2985 => x"0000",
  2986 => x"0000",
  2987 => x"0000",
  2988 => x"0000",
  2989 => x"0000",
  2990 => x"0000",
  2991 => x"0000",
  2992 => x"0000",
  2993 => x"0000",
  2994 => x"0000",
  2995 => x"0000",
  2996 => x"0000",
  2997 => x"0000",
  2998 => x"0000",
  2999 => x"0000",
  3000 => x"0000",
  3001 => x"0000",
  3002 => x"0000",
  3003 => x"0000",
  3004 => x"0000",
  3005 => x"0000",
  3006 => x"0000",
  3007 => x"0000",
  3008 => x"0000",
  3009 => x"0000",
  3010 => x"0000",
  3011 => x"0000",
  3012 => x"0000",
  3013 => x"0000",
  3014 => x"0000",
  3015 => x"0000",
  3016 => x"0000",
  3017 => x"0000",
  3018 => x"0000",
  3019 => x"0000",
  3020 => x"0000",
  3021 => x"0000",
  3022 => x"0000",
  3023 => x"0000",
  3024 => x"0000",
  3025 => x"0000",
  3026 => x"0000",
  3027 => x"0000",
  3028 => x"0000",
  3029 => x"0000",
  3030 => x"0000",
  3031 => x"0000",
  3032 => x"0000",
  3033 => x"0000",
  3034 => x"0000",
  3035 => x"0000",
  3036 => x"0000",
  3037 => x"0000",
  3038 => x"0000",
  3039 => x"0000",
  3040 => x"0000",
  3041 => x"0000",
  3042 => x"0000",
  3043 => x"0000",
  3044 => x"0000",
  3045 => x"0000",
  3046 => x"0000",
  3047 => x"0000",
  3048 => x"0000",
  3049 => x"0000",
  3050 => x"0000",
  3051 => x"0000",
  3052 => x"0000",
  3053 => x"0000",
  3054 => x"0000",
  3055 => x"0000",
  3056 => x"0000",
  3057 => x"0000",
  3058 => x"0000",
  3059 => x"0000",
  3060 => x"0000",
  3061 => x"0000",
  3062 => x"0000",
  3063 => x"0000",
  3064 => x"0000",
  3065 => x"0000",
  3066 => x"0000",
  3067 => x"0000",
  3068 => x"0000",
  3069 => x"0000",
  3070 => x"0000",
  3071 => x"0000",
  3072 => x"0000",
  3073 => x"0000",
  3074 => x"0000",
  3075 => x"0000",
  3076 => x"0000",
  3077 => x"0000",
  3078 => x"0000",
  3079 => x"0000",
  3080 => x"0000",
  3081 => x"0000",
  3082 => x"0000",
  3083 => x"0000",
  3084 => x"0000",
  3085 => x"0000",
  3086 => x"0000",
  3087 => x"0000",
  3088 => x"0000",
  3089 => x"0000",
  3090 => x"0000",
  3091 => x"0000",
  3092 => x"0000",
  3093 => x"0000",
  3094 => x"0000",
  3095 => x"0000",
  3096 => x"0000",
  3097 => x"0000",
  3098 => x"0000",
  3099 => x"0000",
  3100 => x"0000",
  3101 => x"0000",
  3102 => x"0000",
  3103 => x"0000",
  3104 => x"0000",
  3105 => x"0000",
  3106 => x"0000",
  3107 => x"0000",
  3108 => x"0000",
  3109 => x"0000",
  3110 => x"0000",
  3111 => x"0000",
  3112 => x"0000",
  3113 => x"0000",
  3114 => x"0000",
  3115 => x"0000",
  3116 => x"0000",
  3117 => x"0000",
  3118 => x"0000",
  3119 => x"0000",
  3120 => x"0000",
  3121 => x"0000",
  3122 => x"0000",
  3123 => x"0000",
  3124 => x"0000",
  3125 => x"0000",
  3126 => x"0000",
  3127 => x"0000",
  3128 => x"0000",
  3129 => x"0000",
  3130 => x"0000",
  3131 => x"0000",
  3132 => x"0000",
  3133 => x"0000",
  3134 => x"0000",
  3135 => x"0000",
  3136 => x"0000",
  3137 => x"0000",
  3138 => x"0000",
  3139 => x"0000",
  3140 => x"0000",
  3141 => x"0000",
  3142 => x"0000",
  3143 => x"0000",
  3144 => x"0000",
  3145 => x"0000",
  3146 => x"0000",
  3147 => x"0000",
  3148 => x"0000",
  3149 => x"0000",
  3150 => x"0000",
  3151 => x"0000",
  3152 => x"0000",
  3153 => x"0000",
  3154 => x"0000",
  3155 => x"0000",
  3156 => x"0000",
  3157 => x"0000",
  3158 => x"0000",
  3159 => x"0000",
  3160 => x"0000",
  3161 => x"0000",
  3162 => x"0000",
  3163 => x"0000",
  3164 => x"0000",
  3165 => x"0000",
  3166 => x"0000",
  3167 => x"0000",
  3168 => x"0000",
  3169 => x"0000",
  3170 => x"0000",
  3171 => x"0000",
  3172 => x"0000",
  3173 => x"0000",
  3174 => x"0000",
  3175 => x"0000",
  3176 => x"0000",
  3177 => x"0000",
  3178 => x"0000",
  3179 => x"0000",
  3180 => x"0000",
  3181 => x"0000",
  3182 => x"0000",
  3183 => x"0000",
  3184 => x"0000",
  3185 => x"0000",
  3186 => x"0000",
  3187 => x"0000",
  3188 => x"0000",
  3189 => x"0000",
  3190 => x"0000",
  3191 => x"0000",
  3192 => x"0000",
  3193 => x"0000",
  3194 => x"0000",
  3195 => x"0000",
  3196 => x"0000",
  3197 => x"0000",
  3198 => x"0000",
  3199 => x"0000",
  3200 => x"0000",
  3201 => x"0000",
  3202 => x"0000",
  3203 => x"0000",
  3204 => x"0000",
  3205 => x"0000",
  3206 => x"0000",
  3207 => x"0000",
  3208 => x"0000",
  3209 => x"0000",
  3210 => x"0000",
  3211 => x"0000",
  3212 => x"0000",
  3213 => x"0000",
  3214 => x"0000",
  3215 => x"0000",
  3216 => x"0000",
  3217 => x"0000",
  3218 => x"0000",
  3219 => x"0000",
  3220 => x"0000",
  3221 => x"0000",
  3222 => x"0000",
  3223 => x"0000",
  3224 => x"0000",
  3225 => x"0000",
  3226 => x"0000",
  3227 => x"0000",
  3228 => x"0000",
  3229 => x"0000",
  3230 => x"0000",
  3231 => x"0000",
  3232 => x"0000",
  3233 => x"0000",
  3234 => x"0000",
  3235 => x"0000",
  3236 => x"0000",
  3237 => x"0000",
  3238 => x"0000",
  3239 => x"0000",
  3240 => x"0000",
  3241 => x"0000",
  3242 => x"0000",
  3243 => x"0000",
  3244 => x"0000",
  3245 => x"0000",
  3246 => x"0000",
  3247 => x"0000",
  3248 => x"0000",
  3249 => x"0000",
  3250 => x"0000",
  3251 => x"0000",
  3252 => x"0000",
  3253 => x"0000",
  3254 => x"0000",
  3255 => x"0000",
  3256 => x"0000",
  3257 => x"0000",
  3258 => x"0000",
  3259 => x"0000",
  3260 => x"0000",
  3261 => x"0000",
  3262 => x"0000",
  3263 => x"0000",
  3264 => x"0000",
  3265 => x"0000",
  3266 => x"0000",
  3267 => x"0000",
  3268 => x"0000",
  3269 => x"0000",
  3270 => x"0000",
  3271 => x"0000",
  3272 => x"0000",
  3273 => x"0000",
  3274 => x"0000",
  3275 => x"0000",
  3276 => x"0000",
  3277 => x"0000",
  3278 => x"0000",
  3279 => x"0000",
  3280 => x"0000",
  3281 => x"0000",
  3282 => x"0000",
  3283 => x"0000",
  3284 => x"0000",
  3285 => x"0000",
  3286 => x"0000",
  3287 => x"0000",
  3288 => x"0000",
  3289 => x"0000",
  3290 => x"0000",
  3291 => x"0000",
  3292 => x"0000",
  3293 => x"0000",
  3294 => x"0000",
  3295 => x"0000",
  3296 => x"0000",
  3297 => x"0000",
  3298 => x"0000",
  3299 => x"0000",
  3300 => x"0000",
  3301 => x"0000",
  3302 => x"0000",
  3303 => x"0000",
  3304 => x"0000",
  3305 => x"0000",
  3306 => x"0000",
  3307 => x"0000",
  3308 => x"0000",
  3309 => x"0000",
  3310 => x"0000",
  3311 => x"0000",
  3312 => x"0000",
  3313 => x"0000",
  3314 => x"0000",
  3315 => x"0000",
  3316 => x"0000",
  3317 => x"0000",
  3318 => x"0000",
  3319 => x"0000",
  3320 => x"0000",
  3321 => x"0000",
  3322 => x"0000",
  3323 => x"0000",
  3324 => x"0000",
  3325 => x"0000",
  3326 => x"0000",
  3327 => x"0000",
  3328 => x"0000",
  3329 => x"0000",
  3330 => x"0000",
  3331 => x"0000",
  3332 => x"0000",
  3333 => x"0000",
  3334 => x"0000",
  3335 => x"0000",
  3336 => x"0000",
  3337 => x"0000",
  3338 => x"0000",
  3339 => x"0000",
  3340 => x"0000",
  3341 => x"0000",
  3342 => x"0000",
  3343 => x"0000",
  3344 => x"0000",
  3345 => x"0000",
  3346 => x"0000",
  3347 => x"0000",
  3348 => x"0000",
  3349 => x"0000",
  3350 => x"0000",
  3351 => x"0000",
  3352 => x"0000",
  3353 => x"0000",
  3354 => x"0000",
  3355 => x"0000",
  3356 => x"0000",
  3357 => x"0000",
  3358 => x"0000",
  3359 => x"0000",
  3360 => x"0000",
  3361 => x"0000",
  3362 => x"0000",
  3363 => x"0000",
  3364 => x"0000",
  3365 => x"0000",
  3366 => x"0000",
  3367 => x"0000",
  3368 => x"0000",
  3369 => x"0000",
  3370 => x"0000",
  3371 => x"0000",
  3372 => x"0000",
  3373 => x"0000",
  3374 => x"0000",
  3375 => x"0000",
  3376 => x"0000",
  3377 => x"0000",
  3378 => x"0000",
  3379 => x"0000",
  3380 => x"0000",
  3381 => x"0000",
  3382 => x"0000",
  3383 => x"0000",
  3384 => x"0000",
  3385 => x"0000",
  3386 => x"0000",
  3387 => x"0000",
  3388 => x"0000",
  3389 => x"0000",
  3390 => x"0000",
  3391 => x"0000",
  3392 => x"0000",
  3393 => x"0000",
  3394 => x"0000",
  3395 => x"0000",
  3396 => x"0000",
  3397 => x"0000",
  3398 => x"0000",
  3399 => x"0000",
  3400 => x"0000",
  3401 => x"0000",
  3402 => x"0000",
  3403 => x"0000",
  3404 => x"0000",
  3405 => x"0000",
  3406 => x"0000",
  3407 => x"0000",
  3408 => x"0000",
  3409 => x"0000",
  3410 => x"0000",
  3411 => x"0000",
  3412 => x"0000",
  3413 => x"0000",
  3414 => x"0000",
  3415 => x"0000",
  3416 => x"0000",
  3417 => x"0000",
  3418 => x"0000",
  3419 => x"0000",
  3420 => x"0000",
  3421 => x"0000",
  3422 => x"0000",
  3423 => x"0000",
  3424 => x"0000",
  3425 => x"0000",
  3426 => x"0000",
  3427 => x"0000",
  3428 => x"0000",
  3429 => x"0000",
  3430 => x"0000",
  3431 => x"0000",
  3432 => x"0000",
  3433 => x"0000",
  3434 => x"0000",
  3435 => x"0000",
  3436 => x"0000",
  3437 => x"0000",
  3438 => x"0000",
  3439 => x"0000",
  3440 => x"0000",
  3441 => x"0000",
  3442 => x"0000",
  3443 => x"0000",
  3444 => x"0000",
  3445 => x"0000",
  3446 => x"0000",
  3447 => x"0000",
  3448 => x"0000",
  3449 => x"0000",
  3450 => x"0000",
  3451 => x"0000",
  3452 => x"0000",
  3453 => x"0000",
  3454 => x"0000",
  3455 => x"0000",
  3456 => x"0000",
  3457 => x"0000",
  3458 => x"0000",
  3459 => x"0000",
  3460 => x"0000",
  3461 => x"0000",
  3462 => x"0000",
  3463 => x"0000",
  3464 => x"0000",
  3465 => x"0000",
  3466 => x"0000",
  3467 => x"0000",
  3468 => x"0000",
  3469 => x"0000",
  3470 => x"0000",
  3471 => x"0000",
  3472 => x"0000",
  3473 => x"0000",
  3474 => x"0000",
  3475 => x"0000",
  3476 => x"0000",
  3477 => x"0000",
  3478 => x"0000",
  3479 => x"0000",
  3480 => x"0000",
  3481 => x"0000",
  3482 => x"0000",
  3483 => x"0000",
  3484 => x"0000",
  3485 => x"0000",
  3486 => x"0000",
  3487 => x"0000",
  3488 => x"0000",
  3489 => x"0000",
  3490 => x"0000",
  3491 => x"0000",
  3492 => x"0000",
  3493 => x"0000",
  3494 => x"0000",
  3495 => x"0000",
  3496 => x"0000",
  3497 => x"0000",
  3498 => x"0000",
  3499 => x"0000",
  3500 => x"0000",
  3501 => x"0000",
  3502 => x"0000",
  3503 => x"0000",
  3504 => x"0000",
  3505 => x"0000",
  3506 => x"0000",
  3507 => x"0000",
  3508 => x"0000",
  3509 => x"0000",
  3510 => x"0000",
  3511 => x"0000",
  3512 => x"0000",
  3513 => x"0000",
  3514 => x"0000",
  3515 => x"0000",
  3516 => x"0000",
  3517 => x"0000",
  3518 => x"0000",
  3519 => x"0000",
  3520 => x"0000",
  3521 => x"0000",
  3522 => x"0000",
  3523 => x"0000",
  3524 => x"0000",
  3525 => x"0000",
  3526 => x"0000",
  3527 => x"0000",
  3528 => x"0000",
  3529 => x"0000",
  3530 => x"0000",
  3531 => x"0000",
  3532 => x"0000",
  3533 => x"0000",
  3534 => x"0000",
  3535 => x"0000",
  3536 => x"0000",
  3537 => x"0000",
  3538 => x"0000",
  3539 => x"0000",
  3540 => x"0000",
  3541 => x"0000",
  3542 => x"0000",
  3543 => x"0000",
  3544 => x"0000",
  3545 => x"0000",
  3546 => x"0000",
  3547 => x"0000",
  3548 => x"0000",
  3549 => x"0000",
  3550 => x"0000",
  3551 => x"0000",
  3552 => x"0000",
  3553 => x"0000",
  3554 => x"0000",
  3555 => x"0000",
  3556 => x"0000",
  3557 => x"0000",
  3558 => x"0000",
  3559 => x"0000",
  3560 => x"0000",
  3561 => x"0000",
  3562 => x"0000",
  3563 => x"0000",
  3564 => x"0000",
  3565 => x"0000",
  3566 => x"0000",
  3567 => x"0000",
  3568 => x"0000",
  3569 => x"0000",
  3570 => x"0000",
  3571 => x"0000",
  3572 => x"0000",
  3573 => x"0000",
  3574 => x"0000",
  3575 => x"0000",
  3576 => x"0000",
  3577 => x"0000",
  3578 => x"0000",
  3579 => x"0000",
  3580 => x"0000",
  3581 => x"0000",
  3582 => x"0000",
  3583 => x"0000",
  3584 => x"0000",
  3585 => x"0000",
  3586 => x"0000",
  3587 => x"0000",
  3588 => x"0000",
  3589 => x"0000",
  3590 => x"0000",
  3591 => x"0000",
  3592 => x"0000",
  3593 => x"0000",
  3594 => x"0000",
  3595 => x"0000",
  3596 => x"0000",
  3597 => x"0000",
  3598 => x"0000",
  3599 => x"0000",
  3600 => x"0000",
  3601 => x"0000",
  3602 => x"0000",
  3603 => x"0000",
  3604 => x"0000",
  3605 => x"0000",
  3606 => x"0000",
  3607 => x"0000",
  3608 => x"0000",
  3609 => x"0000",
  3610 => x"0000",
  3611 => x"0000",
  3612 => x"0000",
  3613 => x"0000",
  3614 => x"0000",
  3615 => x"0000",
  3616 => x"0000",
  3617 => x"0000",
  3618 => x"0000",
  3619 => x"0000",
  3620 => x"0000",
  3621 => x"0000",
  3622 => x"0000",
  3623 => x"0000",
  3624 => x"0000",
  3625 => x"0000",
  3626 => x"0000",
  3627 => x"0000",
  3628 => x"0000",
  3629 => x"0000",
  3630 => x"0000",
  3631 => x"0000",
  3632 => x"0000",
  3633 => x"0000",
  3634 => x"0000",
  3635 => x"0000",
  3636 => x"0000",
  3637 => x"0000",
  3638 => x"0000",
  3639 => x"0000",
  3640 => x"0000",
  3641 => x"0000",
  3642 => x"0000",
  3643 => x"0000",
  3644 => x"0000",
  3645 => x"0000",
  3646 => x"0000",
  3647 => x"0000",
  3648 => x"0000",
  3649 => x"0000",
  3650 => x"0000",
  3651 => x"0000",
  3652 => x"0000",
  3653 => x"0000",
  3654 => x"0000",
  3655 => x"0000",
  3656 => x"0000",
  3657 => x"0000",
  3658 => x"0000",
  3659 => x"0000",
  3660 => x"0000",
  3661 => x"0000",
  3662 => x"0000",
  3663 => x"0000",
  3664 => x"0000",
  3665 => x"0000",
  3666 => x"0000",
  3667 => x"0000",
  3668 => x"0000",
  3669 => x"0000",
  3670 => x"0000",
  3671 => x"0000",
  3672 => x"0000",
  3673 => x"0000",
  3674 => x"0000",
  3675 => x"0000",
  3676 => x"0000",
  3677 => x"0000",
  3678 => x"0000",
  3679 => x"0000",
  3680 => x"0000",
  3681 => x"0000",
  3682 => x"0000",
  3683 => x"0000",
  3684 => x"0000",
  3685 => x"0000",
  3686 => x"0000",
  3687 => x"0000",
  3688 => x"0000",
  3689 => x"0000",
  3690 => x"0000",
  3691 => x"0000",
  3692 => x"0000",
  3693 => x"0000",
  3694 => x"0000",
  3695 => x"0000",
  3696 => x"0000",
  3697 => x"0000",
  3698 => x"0000",
  3699 => x"0000",
  3700 => x"0000",
  3701 => x"0000",
  3702 => x"0000",
  3703 => x"0000",
  3704 => x"0000",
  3705 => x"0000",
  3706 => x"0000",
  3707 => x"0000",
  3708 => x"0000",
  3709 => x"0000",
  3710 => x"0000",
  3711 => x"0000",
  3712 => x"0000",
  3713 => x"0000",
  3714 => x"0000",
  3715 => x"0000",
  3716 => x"0000",
  3717 => x"0000",
  3718 => x"0000",
  3719 => x"0000",
  3720 => x"0000",
  3721 => x"0000",
  3722 => x"0000",
  3723 => x"0000",
  3724 => x"0000",
  3725 => x"0000",
  3726 => x"0000",
  3727 => x"0000",
  3728 => x"0000",
  3729 => x"0000",
  3730 => x"0000",
  3731 => x"0000",
  3732 => x"0000",
  3733 => x"0000",
  3734 => x"0000",
  3735 => x"0000",
  3736 => x"0000",
  3737 => x"0000",
  3738 => x"0000",
  3739 => x"0000",
  3740 => x"0000",
  3741 => x"0000",
  3742 => x"0000",
  3743 => x"0000",
  3744 => x"0000",
  3745 => x"0000",
  3746 => x"0000",
  3747 => x"0000",
  3748 => x"0000",
  3749 => x"0000",
  3750 => x"0000",
  3751 => x"0000",
  3752 => x"0000",
  3753 => x"0000",
  3754 => x"0000",
  3755 => x"0000",
  3756 => x"0000",
  3757 => x"0000",
  3758 => x"0000",
  3759 => x"0000",
  3760 => x"0000",
  3761 => x"0000",
  3762 => x"0000",
  3763 => x"0000",
  3764 => x"0000",
  3765 => x"0000",
  3766 => x"0000",
  3767 => x"0000",
  3768 => x"0000",
  3769 => x"0000",
  3770 => x"0000",
  3771 => x"0000",
  3772 => x"0000",
  3773 => x"0000",
  3774 => x"0000",
  3775 => x"0000",
  3776 => x"0000",
  3777 => x"0000",
  3778 => x"0000",
  3779 => x"0000",
  3780 => x"0000",
  3781 => x"0000",
  3782 => x"0000",
  3783 => x"0000",
  3784 => x"0000",
  3785 => x"0000",
  3786 => x"0000",
  3787 => x"0000",
  3788 => x"0000",
  3789 => x"0000",
  3790 => x"0000",
  3791 => x"0000",
  3792 => x"0000",
  3793 => x"0000",
  3794 => x"0000",
  3795 => x"0000",
  3796 => x"0000",
  3797 => x"0000",
  3798 => x"0000",
  3799 => x"0000",
  3800 => x"0000",
  3801 => x"0000",
  3802 => x"0000",
  3803 => x"0000",
  3804 => x"0000",
  3805 => x"0000",
  3806 => x"0000",
  3807 => x"0000",
  3808 => x"0000",
  3809 => x"0000",
  3810 => x"0000",
  3811 => x"0000",
  3812 => x"0000",
  3813 => x"0000",
  3814 => x"0000",
  3815 => x"0000",
  3816 => x"0000",
  3817 => x"0000",
  3818 => x"0000",
  3819 => x"0000",
  3820 => x"0000",
  3821 => x"0000",
  3822 => x"0000",
  3823 => x"0000",
  3824 => x"0000",
  3825 => x"0000",
  3826 => x"0000",
  3827 => x"0000",
  3828 => x"0000",
  3829 => x"0000",
  3830 => x"0000",
  3831 => x"0000",
  3832 => x"0000",
  3833 => x"0000",
  3834 => x"0000",
  3835 => x"0000",
  3836 => x"0000",
  3837 => x"0000",
  3838 => x"0000",
  3839 => x"0000",
  3840 => x"0000",
  3841 => x"0000",
  3842 => x"0000",
  3843 => x"0000",
  3844 => x"0000",
  3845 => x"0000",
  3846 => x"0000",
  3847 => x"0000",
  3848 => x"0000",
  3849 => x"0000",
  3850 => x"0000",
  3851 => x"0000",
  3852 => x"0000",
  3853 => x"0000",
  3854 => x"0000",
  3855 => x"0000",
  3856 => x"0000",
  3857 => x"0000",
  3858 => x"0000",
  3859 => x"0000",
  3860 => x"0000",
  3861 => x"0000",
  3862 => x"0000",
  3863 => x"0000",
  3864 => x"0000",
  3865 => x"0000",
  3866 => x"0000",
  3867 => x"0000",
  3868 => x"0000",
  3869 => x"0000",
  3870 => x"0000",
  3871 => x"0000",
  3872 => x"0000",
  3873 => x"0000",
  3874 => x"0000",
  3875 => x"0000",
  3876 => x"0000",
  3877 => x"0000",
  3878 => x"0000",
  3879 => x"0000",
  3880 => x"0000",
  3881 => x"0000",
  3882 => x"0000",
  3883 => x"0000",
  3884 => x"0000",
  3885 => x"0000",
  3886 => x"0000",
  3887 => x"0000",
  3888 => x"0000",
  3889 => x"0000",
  3890 => x"0000",
  3891 => x"0000",
  3892 => x"0000",
  3893 => x"0000",
  3894 => x"0000",
  3895 => x"0000",
  3896 => x"0000",
  3897 => x"0000",
  3898 => x"0000",
  3899 => x"0000",
  3900 => x"0000",
  3901 => x"0000",
  3902 => x"0000",
  3903 => x"0000",
  3904 => x"0000",
  3905 => x"0000",
  3906 => x"0000",
  3907 => x"0000",
  3908 => x"0000",
  3909 => x"0000",
  3910 => x"0000",
  3911 => x"0000",
  3912 => x"0000",
  3913 => x"0000",
  3914 => x"0000",
  3915 => x"0000",
  3916 => x"0000",
  3917 => x"0000",
  3918 => x"0000",
  3919 => x"0000",
  3920 => x"0000",
  3921 => x"0000",
  3922 => x"0000",
  3923 => x"0000",
  3924 => x"0000",
  3925 => x"0000",
  3926 => x"0000",
  3927 => x"0000",
  3928 => x"0000",
  3929 => x"0000",
  3930 => x"0000",
  3931 => x"0000",
  3932 => x"0000",
  3933 => x"0000",
  3934 => x"0000",
  3935 => x"0000",
  3936 => x"0000",
  3937 => x"0000",
  3938 => x"0000",
  3939 => x"0000",
  3940 => x"0000",
  3941 => x"0000",
  3942 => x"0000",
  3943 => x"0000",
  3944 => x"0000",
  3945 => x"0000",
  3946 => x"0000",
  3947 => x"0000",
  3948 => x"0000",
  3949 => x"0000",
  3950 => x"0000",
  3951 => x"0000",
  3952 => x"0000",
  3953 => x"0000",
  3954 => x"0000",
  3955 => x"0000",
  3956 => x"0000",
  3957 => x"0000",
  3958 => x"0000",
  3959 => x"0000",
  3960 => x"0000",
  3961 => x"0000",
  3962 => x"0000",
  3963 => x"0000",
  3964 => x"0000",
  3965 => x"0000",
  3966 => x"0000",
  3967 => x"0000",
  3968 => x"0000",
  3969 => x"0000",
  3970 => x"0000",
  3971 => x"0000",
  3972 => x"0000",
  3973 => x"0000",
  3974 => x"0000",
  3975 => x"0000",
  3976 => x"0000",
  3977 => x"0000",
  3978 => x"0000",
  3979 => x"0000",
  3980 => x"0000",
  3981 => x"0000",
  3982 => x"0000",
  3983 => x"0000",
  3984 => x"0000",
  3985 => x"0000",
  3986 => x"0000",
  3987 => x"0000",
  3988 => x"0000",
  3989 => x"0000",
  3990 => x"0000",
  3991 => x"0000",
  3992 => x"0000",
  3993 => x"0000",
  3994 => x"0000",
  3995 => x"0000",
  3996 => x"0000",
  3997 => x"0000",
  3998 => x"0000",
  3999 => x"0000",
  4000 => x"0000",
  4001 => x"0000",
  4002 => x"0000",
  4003 => x"0000",
  4004 => x"0000",
  4005 => x"0000",
  4006 => x"0000",
  4007 => x"0000",
  4008 => x"0000",
  4009 => x"0000",
  4010 => x"0000",
  4011 => x"0000",
  4012 => x"0000",
  4013 => x"0000",
  4014 => x"0000",
  4015 => x"0000",
  4016 => x"0000",
  4017 => x"0000",
  4018 => x"0000",
  4019 => x"0000",
  4020 => x"0000",
  4021 => x"0000",
  4022 => x"0000",
  4023 => x"0000",
  4024 => x"0000",
  4025 => x"0000",
  4026 => x"0000",
  4027 => x"0000",
  4028 => x"0000",
  4029 => x"0000",
  4030 => x"0000",
  4031 => x"0000",
  4032 => x"0000",
  4033 => x"0000",
  4034 => x"0000",
  4035 => x"0000",
  4036 => x"0000",
  4037 => x"0000",
  4038 => x"0000",
  4039 => x"0000",
  4040 => x"0000",
  4041 => x"0000",
  4042 => x"0000",
  4043 => x"0000",
  4044 => x"0000",
  4045 => x"0000",
  4046 => x"0000",
  4047 => x"0000",
  4048 => x"0000",
  4049 => x"0000",
  4050 => x"0000",
  4051 => x"0000",
  4052 => x"0000",
  4053 => x"0000",
  4054 => x"0000",
  4055 => x"0000",
  4056 => x"0000",
  4057 => x"0000",
  4058 => x"0000",
  4059 => x"0000",
  4060 => x"0000",
  4061 => x"0000",
  4062 => x"0000",
  4063 => x"0000",
  4064 => x"0000",
  4065 => x"0000",
  4066 => x"0000",
  4067 => x"0000",
  4068 => x"0000",
  4069 => x"0000",
  4070 => x"0000",
  4071 => x"0000",
  4072 => x"0000",
  4073 => x"0000",
  4074 => x"0000",
  4075 => x"0000",
  4076 => x"0000",
  4077 => x"0000",
  4078 => x"0000",
  4079 => x"0000",
  4080 => x"0000",
  4081 => x"0000",
  4082 => x"0000",
  4083 => x"0000",
  4084 => x"0000",
  4085 => x"0000",
  4086 => x"0000",
  4087 => x"0000",
  4088 => x"0000",
  4089 => x"0000",
  4090 => x"0000",
  4091 => x"0000",
  4092 => x"0000",
  4093 => x"0000",
  4094 => x"0000",
  4095 => x"0000",
  4096 => x"0000",
  4097 => x"0000",
  4098 => x"0000",
  4099 => x"0000",
  4100 => x"0000",
  4101 => x"0000",
  4102 => x"0000",
  4103 => x"0000",
  4104 => x"0000",
  4105 => x"0000",
  4106 => x"0000",
  4107 => x"0000",
  4108 => x"0000",
  4109 => x"0000",
  4110 => x"0000",
  4111 => x"0000",
  4112 => x"0000",
  4113 => x"0000",
  4114 => x"0000",
  4115 => x"0000",
  4116 => x"0000",
  4117 => x"0000",
  4118 => x"0000",
  4119 => x"0000",
  4120 => x"0000",
  4121 => x"0000",
  4122 => x"0000",
  4123 => x"0000",
  4124 => x"0000",
  4125 => x"0000",
  4126 => x"0000",
  4127 => x"0000",
  4128 => x"0000",
  4129 => x"0000",
  4130 => x"0000",
  4131 => x"0000",
  4132 => x"0000",
  4133 => x"0000",
  4134 => x"0000",
  4135 => x"0000",
  4136 => x"0000",
  4137 => x"0000",
  4138 => x"0000",
  4139 => x"0000",
  4140 => x"0000",
  4141 => x"0000",
  4142 => x"0000",
  4143 => x"0000",
  4144 => x"0000",
  4145 => x"0000",
  4146 => x"0000",
  4147 => x"0000",
  4148 => x"0000",
  4149 => x"0000",
  4150 => x"0000",
  4151 => x"0000",
  4152 => x"0000",
  4153 => x"0000",
  4154 => x"0000",
  4155 => x"0000",
  4156 => x"0000",
  4157 => x"0000",
  4158 => x"0000",
  4159 => x"0000",
  4160 => x"0000",
  4161 => x"0000",
  4162 => x"0000",
  4163 => x"0000",
  4164 => x"0000",
  4165 => x"0000",
  4166 => x"0000",
  4167 => x"0000",
  4168 => x"0000",
  4169 => x"0000",
  4170 => x"0000",
  4171 => x"0000",
  4172 => x"0000",
  4173 => x"0000",
  4174 => x"0000",
  4175 => x"0000",
  4176 => x"0000",
  4177 => x"0000",
  4178 => x"0000",
  4179 => x"0000",
  4180 => x"0000",
  4181 => x"0000",
  4182 => x"0000",
  4183 => x"0000",
  4184 => x"0000",
  4185 => x"0000",
  4186 => x"0000",
  4187 => x"0000",
  4188 => x"0000",
  4189 => x"0000",
  4190 => x"0000",
  4191 => x"0000",
  4192 => x"0000",
  4193 => x"0000",
  4194 => x"0000",
  4195 => x"0000",
  4196 => x"0000",
  4197 => x"0000",
  4198 => x"0000",
  4199 => x"0000",
  4200 => x"0000",
  4201 => x"0000",
  4202 => x"0000",
  4203 => x"0000",
  4204 => x"0000",
  4205 => x"0000",
  4206 => x"0000",
  4207 => x"0000",
  4208 => x"0000",
  4209 => x"0000",
  4210 => x"0000",
  4211 => x"0000",
  4212 => x"0000",
  4213 => x"0000",
  4214 => x"0000",
  4215 => x"0000",
  4216 => x"0000",
  4217 => x"0000",
  4218 => x"0000",
  4219 => x"0000",
  4220 => x"0000",
  4221 => x"0000",
  4222 => x"0000",
  4223 => x"0000",
  4224 => x"0000",
  4225 => x"0000",
  4226 => x"0000",
  4227 => x"0000",
  4228 => x"0000",
  4229 => x"0000",
  4230 => x"0000",
  4231 => x"0000",
  4232 => x"0000",
  4233 => x"0000",
  4234 => x"0000",
  4235 => x"0000",
  4236 => x"0000",
  4237 => x"0000",
  4238 => x"0000",
  4239 => x"0000",
  4240 => x"0000",
  4241 => x"0000",
  4242 => x"0000",
  4243 => x"0000",
  4244 => x"0000",
  4245 => x"0000",
  4246 => x"0000",
  4247 => x"0000",
  4248 => x"0000",
  4249 => x"0000",
  4250 => x"0000",
  4251 => x"0000",
  4252 => x"0000",
  4253 => x"0000",
  4254 => x"0000",
  4255 => x"0000",
  4256 => x"0000",
  4257 => x"0000",
  4258 => x"0000",
  4259 => x"0000",
  4260 => x"0000",
  4261 => x"0000",
  4262 => x"0000",
  4263 => x"0000",
  4264 => x"0000",
  4265 => x"0000",
  4266 => x"0000",
  4267 => x"0000",
  4268 => x"0000",
  4269 => x"0000",
  4270 => x"0000",
  4271 => x"0000",
  4272 => x"0000",
  4273 => x"0000",
  4274 => x"0000",
  4275 => x"0000",
  4276 => x"0000",
  4277 => x"0000",
  4278 => x"0000",
  4279 => x"0000",
  4280 => x"0000",
  4281 => x"0000",
  4282 => x"0000",
  4283 => x"0000",
  4284 => x"0000",
  4285 => x"0000",
  4286 => x"0000",
  4287 => x"0000",
  4288 => x"0000",
  4289 => x"0000",
  4290 => x"0000",
  4291 => x"0000",
  4292 => x"0000",
  4293 => x"0000",
  4294 => x"0000",
  4295 => x"0000",
  4296 => x"0000",
  4297 => x"0000",
  4298 => x"0000",
  4299 => x"0000",
  4300 => x"0000",
  4301 => x"0000",
  4302 => x"0000",
  4303 => x"0000",
  4304 => x"0000",
  4305 => x"0000",
  4306 => x"0000",
  4307 => x"0000",
  4308 => x"0000",
  4309 => x"0000",
  4310 => x"0000",
  4311 => x"0000",
  4312 => x"0000",
  4313 => x"0000",
  4314 => x"0000",
  4315 => x"0000",
  4316 => x"0000",
  4317 => x"0000",
  4318 => x"0000",
  4319 => x"0000",
  4320 => x"0000",
  4321 => x"0000",
  4322 => x"0000",
  4323 => x"0000",
  4324 => x"0000",
  4325 => x"0000",
  4326 => x"0000",
  4327 => x"0000",
  4328 => x"0000",
  4329 => x"0000",
  4330 => x"0000",
  4331 => x"0000",
  4332 => x"0000",
  4333 => x"0000",
  4334 => x"0000",
  4335 => x"0000",
  4336 => x"0000",
  4337 => x"0000",
  4338 => x"0000",
  4339 => x"0000",
  4340 => x"0000",
  4341 => x"0000",
  4342 => x"0000",
  4343 => x"0000",
  4344 => x"0000",
  4345 => x"0000",
  4346 => x"0000",
  4347 => x"0000",
  4348 => x"0000",
  4349 => x"0000",
  4350 => x"0000",
  4351 => x"0000",
  4352 => x"0000",
  4353 => x"0000",
  4354 => x"0000",
  4355 => x"0000",
  4356 => x"0000",
  4357 => x"0000",
  4358 => x"0000",
  4359 => x"0000",
  4360 => x"0000",
  4361 => x"0000",
  4362 => x"0000",
  4363 => x"0000",
  4364 => x"0000",
  4365 => x"0000",
  4366 => x"0000",
  4367 => x"0000",
  4368 => x"0000",
  4369 => x"0000",
  4370 => x"0000",
  4371 => x"0000",
  4372 => x"0000",
  4373 => x"0000",
  4374 => x"0000",
  4375 => x"0000",
  4376 => x"0000",
  4377 => x"0000",
  4378 => x"0000",
  4379 => x"0000",
  4380 => x"0000",
  4381 => x"0000",
  4382 => x"0000",
  4383 => x"0000",
  4384 => x"0000",
  4385 => x"0000",
  4386 => x"0000",
  4387 => x"0000",
  4388 => x"0000",
  4389 => x"0000",
  4390 => x"0000",
  4391 => x"0000",
  4392 => x"0000",
  4393 => x"0000",
  4394 => x"0000",
  4395 => x"0000",
  4396 => x"0000",
  4397 => x"0000",
  4398 => x"0000",
  4399 => x"0000",
  4400 => x"0000",
  4401 => x"0000",
  4402 => x"0000",
  4403 => x"0000",
  4404 => x"0000",
  4405 => x"0000",
  4406 => x"0000",
  4407 => x"0000",
  4408 => x"0000",
  4409 => x"0000",
  4410 => x"0000",
  4411 => x"0000",
  4412 => x"0000",
  4413 => x"0000",
  4414 => x"0000",
  4415 => x"0000",
  4416 => x"0000",
  4417 => x"0000",
  4418 => x"0000",
  4419 => x"0000",
  4420 => x"0000",
  4421 => x"0000",
  4422 => x"0000",
  4423 => x"0000",
  4424 => x"0000",
  4425 => x"0000",
  4426 => x"0000",
  4427 => x"0000",
  4428 => x"0000",
  4429 => x"0000",
  4430 => x"0000",
  4431 => x"0000",
  4432 => x"0000",
  4433 => x"0000",
  4434 => x"0000",
  4435 => x"0000",
  4436 => x"0000",
  4437 => x"0000",
  4438 => x"0000",
  4439 => x"0000",
  4440 => x"0000",
  4441 => x"0000",
  4442 => x"0000",
  4443 => x"0000",
  4444 => x"0000",
  4445 => x"0000",
  4446 => x"0000",
  4447 => x"0000",
  4448 => x"0000",
  4449 => x"0000",
  4450 => x"0000",
  4451 => x"0000",
  4452 => x"0000",
  4453 => x"0000",
  4454 => x"0000",
  4455 => x"0000",
  4456 => x"0000",
  4457 => x"0000",
  4458 => x"0000",
  4459 => x"0000",
  4460 => x"0000",
  4461 => x"0000",
  4462 => x"0000",
  4463 => x"0000",
  4464 => x"0000",
  4465 => x"0000",
  4466 => x"0000",
  4467 => x"0000",
  4468 => x"0000",
  4469 => x"0000",
  4470 => x"0000",
  4471 => x"0000",
  4472 => x"0000",
  4473 => x"0000",
  4474 => x"0000",
  4475 => x"0000",
  4476 => x"0000",
  4477 => x"0000",
  4478 => x"0000",
  4479 => x"0000",
  4480 => x"0000",
  4481 => x"0000",
  4482 => x"0000",
  4483 => x"0000",
  4484 => x"0000",
  4485 => x"0000",
  4486 => x"0000",
  4487 => x"0000",
  4488 => x"0000",
  4489 => x"0000",
  4490 => x"0000",
  4491 => x"0000",
  4492 => x"0000",
  4493 => x"0000",
  4494 => x"0000",
  4495 => x"0000",
  4496 => x"0000",
  4497 => x"0000",
  4498 => x"0000",
  4499 => x"0000",
  4500 => x"0000",
  4501 => x"0000",
  4502 => x"0000",
  4503 => x"0000",
  4504 => x"0000",
  4505 => x"0000",
  4506 => x"0000",
  4507 => x"0000",
  4508 => x"0000",
  4509 => x"0000",
  4510 => x"0000",
  4511 => x"0000",
  4512 => x"0000",
  4513 => x"0000",
  4514 => x"0000",
  4515 => x"0000",
  4516 => x"0000",
  4517 => x"0000",
  4518 => x"0000",
  4519 => x"0000",
  4520 => x"0000",
  4521 => x"0000",
  4522 => x"0000",
  4523 => x"0000",
  4524 => x"0000",
  4525 => x"0000",
  4526 => x"0000",
  4527 => x"0000",
  4528 => x"0000",
  4529 => x"0000",
  4530 => x"0000",
  4531 => x"0000",
  4532 => x"0000",
  4533 => x"0000",
  4534 => x"0000",
  4535 => x"0000",
  4536 => x"0000",
  4537 => x"0000",
  4538 => x"0000",
  4539 => x"0000",
  4540 => x"0000",
  4541 => x"0000",
  4542 => x"0000",
  4543 => x"0000",
  4544 => x"0000",
  4545 => x"0000",
  4546 => x"0000",
  4547 => x"0000",
  4548 => x"0000",
  4549 => x"0000",
  4550 => x"0000",
  4551 => x"0000",
  4552 => x"0000",
  4553 => x"0000",
  4554 => x"0000",
  4555 => x"0000",
  4556 => x"0000",
  4557 => x"0000",
  4558 => x"0000",
  4559 => x"0000",
  4560 => x"0000",
  4561 => x"0000",
  4562 => x"0000",
  4563 => x"0000",
  4564 => x"0000",
  4565 => x"0000",
  4566 => x"0000",
  4567 => x"0000",
  4568 => x"0000",
  4569 => x"0000",
  4570 => x"0000",
  4571 => x"0000",
  4572 => x"0000",
  4573 => x"0000",
  4574 => x"0000",
  4575 => x"0000",
  4576 => x"0000",
  4577 => x"0000",
  4578 => x"0000",
  4579 => x"0000",
  4580 => x"0000",
  4581 => x"0000",
  4582 => x"0000",
  4583 => x"0000",
  4584 => x"0000",
  4585 => x"0000",
  4586 => x"0000",
  4587 => x"0000",
  4588 => x"0000",
  4589 => x"0000",
  4590 => x"0000",
  4591 => x"0000",
  4592 => x"0000",
  4593 => x"0000",
  4594 => x"0000",
  4595 => x"0000",
  4596 => x"0000",
  4597 => x"0000",
  4598 => x"0000",
  4599 => x"0000",
  4600 => x"0000",
  4601 => x"0000",
  4602 => x"0000",
  4603 => x"0000",
  4604 => x"0000",
  4605 => x"0000",
  4606 => x"0000",
  4607 => x"0000",
  4608 => x"0000",
  4609 => x"0000",
  4610 => x"0000",
  4611 => x"0000",
  4612 => x"0000",
  4613 => x"0000",
  4614 => x"0000",
  4615 => x"0000",
  4616 => x"0000",
  4617 => x"0000",
  4618 => x"0000",
  4619 => x"0000",
  4620 => x"0000",
  4621 => x"0000",
  4622 => x"0000",
  4623 => x"0000",
  4624 => x"0000",
  4625 => x"0000",
  4626 => x"0000",
  4627 => x"0000",
  4628 => x"0000",
  4629 => x"0000",
  4630 => x"0000",
  4631 => x"0000",
  4632 => x"0000",
  4633 => x"0000",
  4634 => x"0000",
  4635 => x"0000",
  4636 => x"0000",
  4637 => x"0000",
  4638 => x"0000",
  4639 => x"0000",
  4640 => x"0000",
  4641 => x"0000",
  4642 => x"0000",
  4643 => x"0000",
  4644 => x"0000",
  4645 => x"0000",
  4646 => x"0000",
  4647 => x"0000",
  4648 => x"0000",
  4649 => x"0000",
  4650 => x"0000",
  4651 => x"0000",
  4652 => x"0000",
  4653 => x"0000",
  4654 => x"0000",
  4655 => x"0000",
  4656 => x"0000",
  4657 => x"0000",
  4658 => x"0000",
  4659 => x"0000",
  4660 => x"0000",
  4661 => x"0000",
  4662 => x"0000",
  4663 => x"0000",
  4664 => x"0000",
  4665 => x"0000",
  4666 => x"0000",
  4667 => x"0000",
  4668 => x"0000",
  4669 => x"0000",
  4670 => x"0000",
  4671 => x"0000",
  4672 => x"0000",
  4673 => x"0000",
  4674 => x"0000",
  4675 => x"0000",
  4676 => x"0000",
  4677 => x"0000",
  4678 => x"0000",
  4679 => x"0000",
  4680 => x"0000",
  4681 => x"0000",
  4682 => x"0000",
  4683 => x"0000",
  4684 => x"0000",
  4685 => x"0000",
  4686 => x"0000",
  4687 => x"0000",
  4688 => x"0000",
  4689 => x"0000",
  4690 => x"0000",
  4691 => x"0000",
  4692 => x"0000",
  4693 => x"0000",
  4694 => x"0000",
  4695 => x"0000",
  4696 => x"0000",
  4697 => x"0000",
  4698 => x"0000",
  4699 => x"0000",
  4700 => x"0000",
  4701 => x"0000",
  4702 => x"0000",
  4703 => x"0000",
  4704 => x"0000",
  4705 => x"0000",
  4706 => x"0000",
  4707 => x"0000",
  4708 => x"0000",
  4709 => x"0000",
  4710 => x"0000",
  4711 => x"0000",
  4712 => x"0000",
  4713 => x"0000",
  4714 => x"0000",
  4715 => x"0000",
  4716 => x"0000",
  4717 => x"0000",
  4718 => x"0000",
  4719 => x"0000",
  4720 => x"0000",
  4721 => x"0000",
  4722 => x"0000",
  4723 => x"0000",
  4724 => x"0000",
  4725 => x"0000",
  4726 => x"0000",
  4727 => x"0000",
  4728 => x"0000",
  4729 => x"0000",
  4730 => x"0000",
  4731 => x"0000",
  4732 => x"0000",
  4733 => x"0000",
  4734 => x"0000",
  4735 => x"0000",
  4736 => x"0000",
  4737 => x"0000",
  4738 => x"0000",
  4739 => x"0000",
  4740 => x"0000",
  4741 => x"0000",
  4742 => x"0000",
  4743 => x"0000",
  4744 => x"0000",
  4745 => x"0000",
  4746 => x"0000",
  4747 => x"0000",
  4748 => x"0000",
  4749 => x"0000",
  4750 => x"0000",
  4751 => x"0000",
  4752 => x"0000",
  4753 => x"0000",
  4754 => x"0000",
  4755 => x"0000",
  4756 => x"0000",
  4757 => x"0000",
  4758 => x"0000",
  4759 => x"0000",
  4760 => x"0000",
  4761 => x"0000",
  4762 => x"0000",
  4763 => x"0000",
  4764 => x"0000",
  4765 => x"0000",
  4766 => x"0000",
  4767 => x"0000",
  4768 => x"0000",
  4769 => x"0000",
  4770 => x"0000",
  4771 => x"0000",
  4772 => x"0000",
  4773 => x"0000",
  4774 => x"0000",
  4775 => x"0000",
  4776 => x"0000",
  4777 => x"0000",
  4778 => x"0000",
  4779 => x"0000",
  4780 => x"0000",
  4781 => x"0000",
  4782 => x"0000",
  4783 => x"0000",
  4784 => x"0000",
  4785 => x"0000",
  4786 => x"0000",
  4787 => x"0000",
  4788 => x"0000",
  4789 => x"0000",
  4790 => x"0000",
  4791 => x"0000",
  4792 => x"0000",
  4793 => x"0000",
  4794 => x"0000",
  4795 => x"0000",
  4796 => x"0000",
  4797 => x"0000",
  4798 => x"0000",
  4799 => x"0000",
  4800 => x"0000",
  4801 => x"0000",
  4802 => x"0000",
  4803 => x"0000",
  4804 => x"0050",
  4805 => x"0000",
  4806 => x"8870",
  4807 => x"0000",
  4808 => x"0050",
  4809 => x"0000",
  4810 => x"7088",
  4811 => x"0000",
  4812 => x"50F8",
  4813 => x"F8F8",
  4814 => x"F870",
  4815 => x"2000",
  4816 => x"2070",
  4817 => x"F8F8",
  4818 => x"F870",
  4819 => x"2000",
  4820 => x"7070",
  4821 => x"20F8",
  4822 => x"F820",
  4823 => x"7000",
  4824 => x"2070",
  4825 => x"F8F8",
  4826 => x"7020",
  4827 => x"7000",
  4828 => x"0000",
  4829 => x"7070",
  4830 => x"7000",
  4831 => x"0000",
  4832 => x"F8F8",
  4833 => x"8888",
  4834 => x"88F8",
  4835 => x"F800",
  4836 => x"0000",
  4837 => x"7050",
  4838 => x"7000",
  4839 => x"0000",
  4840 => x"F8F8",
  4841 => x"88A8",
  4842 => x"88F8",
  4843 => x"F800",
  4844 => x"2070",
  4845 => x"A820",
  4846 => x"7088",
  4847 => x"7000",
  4848 => x"7088",
  4849 => x"7020",
  4850 => x"20F8",
  4851 => x"2000",
  4852 => x"3838",
  4853 => x"2020",
  4854 => x"60E0",
  4855 => x"6000",
  4856 => x"7878",
  4857 => x"4858",
  4858 => x"58C0",
  4859 => x"C000",
  4860 => x"00A8",
  4861 => x"5088",
  4862 => x"50A8",
  4863 => x"0000",
  4864 => x"4060",
  4865 => x"7078",
  4866 => x"7060",
  4867 => x"4000",
  4868 => x"1030",
  4869 => x"70F0",
  4870 => x"7030",
  4871 => x"1000",
  4872 => x"2070",
  4873 => x"A820",
  4874 => x"A870",
  4875 => x"2000",
  4876 => x"5050",
  4877 => x"5050",
  4878 => x"0050",
  4879 => x"5000",
  4880 => x"78E8",
  4881 => x"E878",
  4882 => x"2828",
  4883 => x"2800",
  4884 => x"78C8",
  4885 => x"A050",
  4886 => x"2898",
  4887 => x"F000",
  4888 => x"0000",
  4889 => x"0000",
  4890 => x"F8F8",
  4891 => x"F800",
  4892 => x"2070",
  4893 => x"2020",
  4894 => x"7020",
  4895 => x"F800",
  4896 => x"2070",
  4897 => x"F820",
  4898 => x"2020",
  4899 => x"2000",
  4900 => x"2020",
  4901 => x"2020",
  4902 => x"F870",
  4903 => x"2000",
  4904 => x"0020",
  4905 => x"30F8",
  4906 => x"3020",
  4907 => x"0000",
  4908 => x"0020",
  4909 => x"60F8",
  4910 => x"6020",
  4911 => x"0000",
  4912 => x"0000",
  4913 => x"4078",
  4914 => x"0000",
  4915 => x"0000",
  4916 => x"0000",
  4917 => x"50F8",
  4918 => x"5000",
  4919 => x"0000",
  4920 => x"0020",
  4921 => x"2070",
  4922 => x"70F8",
  4923 => x"F800",
  4924 => x"F8F8",
  4925 => x"7070",
  4926 => x"2020",
  4927 => x"0000",
  4928 => x"0000",
  4929 => x"0000",
  4930 => x"0000",
  4931 => x"0000",
  4932 => x"1818",
  4933 => x"1818",
  4934 => x"0000",
  4935 => x"1800",
  4936 => x"6666",
  4937 => x"6600",
  4938 => x"0000",
  4939 => x"0000",
  4940 => x"6666",
  4941 => x"FF66",
  4942 => x"FF66",
  4943 => x"6600",
  4944 => x"183E",
  4945 => x"603C",
  4946 => x"067C",
  4947 => x"1800",
  4948 => x"6266",
  4949 => x"0C18",
  4950 => x"3066",
  4951 => x"4600",
  4952 => x"3C66",
  4953 => x"3C38",
  4954 => x"6766",
  4955 => x"3F00",
  4956 => x"060C",
  4957 => x"1800",
  4958 => x"0000",
  4959 => x"0000",
  4960 => x"0C18",
  4961 => x"3030",
  4962 => x"3018",
  4963 => x"0C00",
  4964 => x"3018",
  4965 => x"0C0C",
  4966 => x"0C18",
  4967 => x"3000",
  4968 => x"0066",
  4969 => x"3CFF",
  4970 => x"3C66",
  4971 => x"0000",
  4972 => x"0018",
  4973 => x"187E",
  4974 => x"1818",
  4975 => x"0000",
  4976 => x"0000",
  4977 => x"0000",
  4978 => x"0018",
  4979 => x"1830",
  4980 => x"0000",
  4981 => x"007E",
  4982 => x"0000",
  4983 => x"0000",
  4984 => x"0000",
  4985 => x"0000",
  4986 => x"0018",
  4987 => x"1800",
  4988 => x"0003",
  4989 => x"060C",
  4990 => x"1830",
  4991 => x"6000",
  4992 => x"3C66",
  4993 => x"6E76",
  4994 => x"6666",
  4995 => x"3C00",
  4996 => x"1818",
  4997 => x"3818",
  4998 => x"1818",
  4999 => x"7E00",
  5000 => x"3C66",
  5001 => x"060C",
  5002 => x"3060",
  5003 => x"7E00",
  5004 => x"3C66",
  5005 => x"061C",
  5006 => x"0666",
  5007 => x"3C00",
  5008 => x"060E",
  5009 => x"1E66",
  5010 => x"7F06",
  5011 => x"0600",
  5012 => x"7E60",
  5013 => x"7C06",
  5014 => x"0666",
  5015 => x"3C00",
  5016 => x"3C66",
  5017 => x"607C",
  5018 => x"6666",
  5019 => x"3C00",
  5020 => x"7E66",
  5021 => x"0C18",
  5022 => x"1818",
  5023 => x"1800",
  5024 => x"3C66",
  5025 => x"663C",
  5026 => x"6666",
  5027 => x"3C00",
  5028 => x"3C66",
  5029 => x"663E",
  5030 => x"0666",
  5031 => x"3C00",
  5032 => x"0000",
  5033 => x"1800",
  5034 => x"0018",
  5035 => x"0000",
  5036 => x"0000",
  5037 => x"1800",
  5038 => x"0018",
  5039 => x"1830",
  5040 => x"0E18",
  5041 => x"3060",
  5042 => x"3018",
  5043 => x"0E00",
  5044 => x"0000",
  5045 => x"7E00",
  5046 => x"7E00",
  5047 => x"0000",
  5048 => x"7018",
  5049 => x"0C06",
  5050 => x"0C18",
  5051 => x"7000",
  5052 => x"3C66",
  5053 => x"060C",
  5054 => x"1800",
  5055 => x"1800",
  5056 => x"3C66",
  5057 => x"6E6E",
  5058 => x"6062",
  5059 => x"3C00",
  5060 => x"183C",
  5061 => x"667E",
  5062 => x"6666",
  5063 => x"6600",
  5064 => x"7C66",
  5065 => x"667C",
  5066 => x"6666",
  5067 => x"7C00",
  5068 => x"3C66",
  5069 => x"6060",
  5070 => x"6066",
  5071 => x"3C00",
  5072 => x"786C",
  5073 => x"6666",
  5074 => x"666C",
  5075 => x"7800",
  5076 => x"7E60",
  5077 => x"6078",
  5078 => x"6060",
  5079 => x"7E00",
  5080 => x"7E60",
  5081 => x"6078",
  5082 => x"6060",
  5083 => x"6000",
  5084 => x"3C66",
  5085 => x"606E",
  5086 => x"6666",
  5087 => x"3C00",
  5088 => x"6666",
  5089 => x"667E",
  5090 => x"6666",
  5091 => x"6600",
  5092 => x"3C18",
  5093 => x"1818",
  5094 => x"1818",
  5095 => x"3C00",
  5096 => x"1E0C",
  5097 => x"0C0C",
  5098 => x"0C6C",
  5099 => x"3800",
  5100 => x"666C",
  5101 => x"7870",
  5102 => x"786C",
  5103 => x"6600",
  5104 => x"6060",
  5105 => x"6060",
  5106 => x"6060",
  5107 => x"7E00",
  5108 => x"6377",
  5109 => x"7F6B",
  5110 => x"6363",
  5111 => x"6300",
  5112 => x"6676",
  5113 => x"7E7E",
  5114 => x"6E66",
  5115 => x"6600",
  5116 => x"3C66",
  5117 => x"6666",
  5118 => x"6666",
  5119 => x"3C00",
  5120 => x"7C66",
  5121 => x"667C",
  5122 => x"6060",
  5123 => x"6000",
  5124 => x"3C66",
  5125 => x"6666",
  5126 => x"663C",
  5127 => x"0E00",
  5128 => x"7C66",
  5129 => x"667C",
  5130 => x"786C",
  5131 => x"6600",
  5132 => x"3C66",
  5133 => x"603C",
  5134 => x"0666",
  5135 => x"3C00",
  5136 => x"7E18",
  5137 => x"1818",
  5138 => x"1818",
  5139 => x"1800",
  5140 => x"6666",
  5141 => x"6666",
  5142 => x"6666",
  5143 => x"3C00",
  5144 => x"6666",
  5145 => x"6666",
  5146 => x"663C",
  5147 => x"1800",
  5148 => x"6363",
  5149 => x"636B",
  5150 => x"7F77",
  5151 => x"6300",
  5152 => x"6666",
  5153 => x"3C18",
  5154 => x"3C66",
  5155 => x"6600",
  5156 => x"6666",
  5157 => x"663C",
  5158 => x"1818",
  5159 => x"1800",
  5160 => x"7E06",
  5161 => x"0C18",
  5162 => x"3060",
  5163 => x"7E00",
  5164 => x"3C30",
  5165 => x"3030",
  5166 => x"3030",
  5167 => x"3C00",
  5168 => x"0060",
  5169 => x"3018",
  5170 => x"0C06",
  5171 => x"0300",
  5172 => x"3C0C",
  5173 => x"0C0C",
  5174 => x"0C0C",
  5175 => x"3C00",
  5176 => x"0018",
  5177 => x"3C7E",
  5178 => x"1818",
  5179 => x"1818",
  5180 => x"0000",
  5181 => x"0000",
  5182 => x"0000",
  5183 => x"00FF",
  5184 => x"6030",
  5185 => x"1800",
  5186 => x"0000",
  5187 => x"0000",
  5188 => x"0000",
  5189 => x"3C06",
  5190 => x"3E66",
  5191 => x"3E00",
  5192 => x"0060",
  5193 => x"607C",
  5194 => x"6666",
  5195 => x"7C00",
  5196 => x"0000",
  5197 => x"3C60",
  5198 => x"6060",
  5199 => x"3C00",
  5200 => x"0006",
  5201 => x"063E",
  5202 => x"6666",
  5203 => x"3E00",
  5204 => x"0000",
  5205 => x"3C66",
  5206 => x"7E60",
  5207 => x"3C00",
  5208 => x"000E",
  5209 => x"183E",
  5210 => x"1818",
  5211 => x"1800",
  5212 => x"0000",
  5213 => x"3E66",
  5214 => x"663E",
  5215 => x"067C",
  5216 => x"0060",
  5217 => x"607C",
  5218 => x"6666",
  5219 => x"6600",
  5220 => x"0018",
  5221 => x"0038",
  5222 => x"1818",
  5223 => x"3C00",
  5224 => x"0006",
  5225 => x"0006",
  5226 => x"0606",
  5227 => x"063C",
  5228 => x"0060",
  5229 => x"606C",
  5230 => x"786C",
  5231 => x"6600",
  5232 => x"0038",
  5233 => x"1818",
  5234 => x"1818",
  5235 => x"3C00",
  5236 => x"0000",
  5237 => x"667F",
  5238 => x"7F6B",
  5239 => x"6300",
  5240 => x"0000",
  5241 => x"7C66",
  5242 => x"6666",
  5243 => x"6600",
  5244 => x"0000",
  5245 => x"3C66",
  5246 => x"6666",
  5247 => x"3C00",
  5248 => x"0000",
  5249 => x"7C66",
  5250 => x"667C",
  5251 => x"6060",
  5252 => x"0000",
  5253 => x"3E66",
  5254 => x"663E",
  5255 => x"0606",
  5256 => x"0000",
  5257 => x"7C66",
  5258 => x"6060",
  5259 => x"6000",
  5260 => x"0000",
  5261 => x"3E60",
  5262 => x"3C06",
  5263 => x"7C00",
  5264 => x"0018",
  5265 => x"7E18",
  5266 => x"1818",
  5267 => x"0E00",
  5268 => x"0000",
  5269 => x"6666",
  5270 => x"6666",
  5271 => x"3E00",
  5272 => x"0000",
  5273 => x"6666",
  5274 => x"663C",
  5275 => x"1800",
  5276 => x"0000",
  5277 => x"636B",
  5278 => x"7F3E",
  5279 => x"3600",
  5280 => x"0000",
  5281 => x"663C",
  5282 => x"183C",
  5283 => x"6600",
  5284 => x"0000",
  5285 => x"6666",
  5286 => x"663E",
  5287 => x"0C78",
  5288 => x"0000",
  5289 => x"7E0C",
  5290 => x"1830",
  5291 => x"7E00",
  5292 => x"1C30",
  5293 => x"3060",
  5294 => x"3030",
  5295 => x"1C00",
  5296 => x"1818",
  5297 => x"1818",
  5298 => x"1818",
  5299 => x"1818",
  5300 => x"380C",
  5301 => x"0C06",
  5302 => x"0C0C",
  5303 => x"3800",
  5304 => x"0032",
  5305 => x"4C00",
  5306 => x"0000",
  5307 => x"0000",
  5308 => x"0020",
  5309 => x"5088",
  5310 => x"8888",
  5311 => x"F800",
  5312 => x"7088",
  5313 => x"8088",
  5314 => x"7020",
  5315 => x"C000",
  5316 => x"0070",
  5317 => x"8088",
  5318 => x"7020",
  5319 => x"C000",
  5320 => x"1448",
  5321 => x"88C8",
  5322 => x"A898",
  5323 => x"8800",
  5324 => x"2850",
  5325 => x"00B0",
  5326 => x"C888",
  5327 => x"8800",
  5328 => x"1020",
  5329 => x"7088",
  5330 => x"F888",
  5331 => x"8800",
  5332 => x"4020",
  5333 => x"7088",
  5334 => x"F888",
  5335 => x"8800",
  5336 => x"5000",
  5337 => x"7088",
  5338 => x"F888",
  5339 => x"8800",
  5340 => x"2050",
  5341 => x"0070",
  5342 => x"88F8",
  5343 => x"8800",
  5344 => x"1020",
  5345 => x"F880",
  5346 => x"F080",
  5347 => x"F800",
  5348 => x"4020",
  5349 => x"F880",
  5350 => x"F080",
  5351 => x"F800",
  5352 => x"5000",
  5353 => x"F880",
  5354 => x"F080",
  5355 => x"F800",
  5356 => x"2050",
  5357 => x"F880",
  5358 => x"F080",
  5359 => x"F800",
  5360 => x"1020",
  5361 => x"F820",
  5362 => x"2020",
  5363 => x"F800",
  5364 => x"4020",
  5365 => x"F820",
  5366 => x"2020",
  5367 => x"F800",
  5368 => x"5000",
  5369 => x"F820",
  5370 => x"2020",
  5371 => x"F800",
  5372 => x"2050",
  5373 => x"F820",
  5374 => x"2020",
  5375 => x"F800",
  5376 => x"1020",
  5377 => x"7088",
  5378 => x"8888",
  5379 => x"7000",
  5380 => x"4020",
  5381 => x"7088",
  5382 => x"8888",
  5383 => x"7000",
  5384 => x"5000",
  5385 => x"7088",
  5386 => x"8888",
  5387 => x"7000",
  5388 => x"2050",
  5389 => x"7088",
  5390 => x"8888",
  5391 => x"7000",
  5392 => x"1020",
  5393 => x"8888",
  5394 => x"8888",
  5395 => x"7000",
  5396 => x"4020",
  5397 => x"8888",
  5398 => x"8888",
  5399 => x"7000",
  5400 => x"5000",
  5401 => x"8888",
  5402 => x"8888",
  5403 => x"7000",
  5404 => x"2050",
  5405 => x"0088",
  5406 => x"8888",
  5407 => x"7000",
  5408 => x"1020",
  5409 => x"7008",
  5410 => x"7888",
  5411 => x"7800",
  5412 => x"4020",
  5413 => x"7008",
  5414 => x"7888",
  5415 => x"7800",
  5416 => x"5000",
  5417 => x"7008",
  5418 => x"7888",
  5419 => x"7800",
  5420 => x"2050",
  5421 => x"7008",
  5422 => x"7888",
  5423 => x"7800",
  5424 => x"1020",
  5425 => x"7884",
  5426 => x"FC80",
  5427 => x"7C00",
  5428 => x"2010",
  5429 => x"7884",
  5430 => x"FC80",
  5431 => x"7C00",
  5432 => x"5000",
  5433 => x"7884",
  5434 => x"FC80",
  5435 => x"7C00",
  5436 => x"2050",
  5437 => x"7884",
  5438 => x"FC80",
  5439 => x"7C00",
  5440 => x"1020",
  5441 => x"0060",
  5442 => x"2020",
  5443 => x"7000",
  5444 => x"4020",
  5445 => x"0060",
  5446 => x"2020",
  5447 => x"7000",
  5448 => x"0050",
  5449 => x"0060",
  5450 => x"2020",
  5451 => x"7000",
  5452 => x"2050",
  5453 => x"0060",
  5454 => x"2020",
  5455 => x"7000",
  5456 => x"1020",
  5457 => x"0070",
  5458 => x"8888",
  5459 => x"7000",
  5460 => x"4020",
  5461 => x"0070",
  5462 => x"8888",
  5463 => x"7000",
  5464 => x"0050",
  5465 => x"0070",
  5466 => x"8888",
  5467 => x"7000",
  5468 => x"2050",
  5469 => x"0070",
  5470 => x"8888",
  5471 => x"7000",
  5472 => x"1020",
  5473 => x"0088",
  5474 => x"8898",
  5475 => x"6800",
  5476 => x"4020",
  5477 => x"0088",
  5478 => x"8898",
  5479 => x"6800",
  5480 => x"0050",
  5481 => x"0088",
  5482 => x"8898",
  5483 => x"6800",
  5484 => x"2050",
  5485 => x"0088",
  5486 => x"8898",
  5487 => x"6800",
  5488 => x"5000",
  5489 => x"8850",
  5490 => x"2020",
  5491 => x"2000",
  5492 => x"5000",
  5493 => x"8850",
  5494 => x"2040",
  5495 => x"8000",
  5496 => x"2000",
  5497 => x"2040",
  5498 => x"8088",
  5499 => x"7000",
  5500 => x"2020",
  5501 => x"0020",
  5502 => x"2020",
  5503 => x"2000",
  5504 => x"0000",
  5505 => x"4890",
  5506 => x"4800",
  5507 => x"0000",
  5508 => x"0000",
  5509 => x"9048",
  5510 => x"9000",
  5511 => x"0000",
  5512 => x"8822",
  5513 => x"8822",
  5514 => x"8822",
  5515 => x"8822",
  5516 => x"AA55",
  5517 => x"AA55",
  5518 => x"AA55",
  5519 => x"AA54",
  5520 => x"CCFF",
  5521 => x"33CC",
  5522 => x"FF33",
  5523 => x"CCFF",
  5524 => x"3030",
  5525 => x"3030",
  5526 => x"3030",
  5527 => x"3030",
  5528 => x"0000",
  5529 => x"00FC",
  5530 => x"FC00",
  5531 => x"0000",
  5532 => x"3030",
  5533 => x"303C",
  5534 => x"3C00",
  5535 => x"0000",
  5536 => x"3030",
  5537 => x"30F0",
  5538 => x"F000",
  5539 => x"0000",
  5540 => x"0000",
  5541 => x"003C",
  5542 => x"3C30",
  5543 => x"3030",
  5544 => x"0000",
  5545 => x"00F0",
  5546 => x"F030",
  5547 => x"3030",
  5548 => x"3030",
  5549 => x"30F0",
  5550 => x"F030",
  5551 => x"3030",
  5552 => x"3030",
  5553 => x"30FC",
  5554 => x"FC00",
  5555 => x"0000",
  5556 => x"3030",
  5557 => x"303C",
  5558 => x"3C30",
  5559 => x"3030",
  5560 => x"0000",
  5561 => x"00FC",
  5562 => x"FC30",
  5563 => x"3030",
  5564 => x"3030",
  5565 => x"30FC",
  5566 => x"FC30",
  5567 => x"3030",
  5568 => x"3030",
  5569 => x"3030",
  5570 => x"3000",
  5571 => x"0000",
  5572 => x"0000",
  5573 => x"00F0",
  5574 => x"F000",
  5575 => x"0000",
  5576 => x"0000",
  5577 => x"003C",
  5578 => x"3C00",
  5579 => x"0000",
  5580 => x"0000",
  5581 => x"0030",
  5582 => x"3030",
  5583 => x"3030",
  5584 => x"FC84",
  5585 => x"8484",
  5586 => x"8484",
  5587 => x"84FC",
  5588 => x"FCFC",
  5589 => x"CCCC",
  5590 => x"CCCC",
  5591 => x"FCFC",
  5592 => x"FCFC",
  5593 => x"FCFC",
  5594 => x"FCFC",
  5595 => x"FCFC",
  5596 => x"FCFC",
  5597 => x"FCFC",
  5598 => x"0000",
  5599 => x"0000",
  5600 => x"E0E0",
  5601 => x"E0E0",
  5602 => x"E0E0",
  5603 => x"E0E0",
  5604 => x"1C1C",
  5605 => x"1C1C",
  5606 => x"1C1C",
  5607 => x"1C1C",
  5608 => x"0000",
  5609 => x"0000",
  5610 => x"FCFC",
  5611 => x"FCFC",
  5612 => x"0000",
  5613 => x"6890",
  5614 => x"9090",
  5615 => x"6800",
  5616 => x"3048",
  5617 => x"4870",
  5618 => x"4868",
  5619 => x"5000",
  5620 => x"00F8",
  5621 => x"8080",
  5622 => x"8080",
  5623 => x"8000",
  5624 => x"0040",
  5625 => x"A810",
  5626 => x"1010",
  5627 => x"1000",
  5628 => x"2020",
  5629 => x"5050",
  5630 => x"8888",
  5631 => x"F800",
  5632 => x"7088",
  5633 => x"6010",
  5634 => x"7088",
  5635 => x"7000",
  5636 => x"0000",
  5637 => x"7880",
  5638 => x"F880",
  5639 => x"7800",
  5640 => x"2018",
  5641 => x"2040",
  5642 => x"3008",
  5643 => x"7000",
  5644 => x"7088",
  5645 => x"88F8",
  5646 => x"8888",
  5647 => x"7000",
  5648 => x"0000",
  5649 => x"C040",
  5650 => x"4050",
  5651 => x"2000",
  5652 => x"2020",
  5653 => x"5050",
  5654 => x"8888",
  5655 => x"8800",
  5656 => x"00C0",
  5657 => x"2020",
  5658 => x"5048",
  5659 => x"8800",
  5660 => x"0000",
  5661 => x"9080",
  5662 => x"90F8",
  5663 => x"8000",
  5664 => x"00F8",
  5665 => x"8888",
  5666 => x"8888",
  5667 => x"8800",
  5668 => x"0000",
  5669 => x"00F8",
  5670 => x"5050",
  5671 => x"5000",
  5672 => x"FC40",
  5673 => x"2010",
  5674 => x"2040",
  5675 => x"F800",
  5676 => x"0000",
  5677 => x"7890",
  5678 => x"9090",
  5679 => x"6000",
  5680 => x"0000",
  5681 => x"78A0",
  5682 => x"2020",
  5683 => x"1800",
  5684 => x"2020",
  5685 => x"70A8",
  5686 => x"7020",
  5687 => x"2000",
  5688 => x"8048",
  5689 => x"5020",
  5690 => x"5090",
  5691 => x"0800",
  5692 => x"0070",
  5693 => x"8888",
  5694 => x"8850",
  5695 => x"D800",
  5696 => x"00F8",
  5697 => x"00F8",
  5698 => x"00F8",
  5699 => x"0000",
  5700 => x"0020",
  5701 => x"20F8",
  5702 => x"2020",
  5703 => x"F800",
  5704 => x"C030",
  5705 => x"0830",
  5706 => x"C000",
  5707 => x"F800",
  5708 => x"1860",
  5709 => x"8060",
  5710 => x"1800",
  5711 => x"F800",
  5712 => x"0020",
  5713 => x"00F8",
  5714 => x"0020",
  5715 => x"0000",
  5716 => x"3048",
  5717 => x"3000",
  5718 => x"0000",
  5719 => x"0000",
  5720 => x"0018",
  5721 => x"1010",
  5722 => x"9050",
  5723 => x"2000",
  5724 => x"6010",
  5725 => x"2070",
  5726 => x"0000",
  5727 => x"0000",
  5728 => x"7088",
  5729 => x"8890",
  5730 => x"8888",
  5731 => x"88B0",
  5732 => x"0020",
  5733 => x"70A0",
  5734 => x"A070",
  5735 => x"2000",
  5736 => x"3C50",
  5737 => x"90FC",
  5738 => x"9090",
  5739 => x"9C00",
  5740 => x"7C90",
  5741 => x"909C",
  5742 => x"9090",
  5743 => x"7C00",
  5744 => x"7088",
  5745 => x"80F0",
  5746 => x"4040",
  5747 => x"F800",
  5748 => x"8888",
  5749 => x"50F8",
  5750 => x"20F8",
  5751 => x"2000",
  5752 => x"1028",
  5753 => x"2020",
  5754 => x"20A0",
  5755 => x"4000",
  5756 => x"F880",
  5757 => x"80F0",
  5758 => x"8888",
  5759 => x"F000",
  5760 => x"F050",
  5761 => x"5090",
  5762 => x"90F8",
  5763 => x"8800",
  5764 => x"A8A8",
  5765 => x"70A8",
  5766 => x"A8A8",
  5767 => x"A800",
  5768 => x"7088",
  5769 => x"0830",
  5770 => x"0888",
  5771 => x"7000",
  5772 => x"8888",
  5773 => x"C8A8",
  5774 => x"9888",
  5775 => x"8800",
  5776 => x"5020",
  5777 => x"88C8",
  5778 => x"A898",
  5779 => x"8800",
  5780 => x"7848",
  5781 => x"4848",
  5782 => x"4848",
  5783 => x"C800",
  5784 => x"8888",
  5785 => x"8888",
  5786 => x"88F8",
  5787 => x"0800",
  5788 => x"8888",
  5789 => x"8878",
  5790 => x"0808",
  5791 => x"0800",
  5792 => x"A8A8",
  5793 => x"A8A8",
  5794 => x"A8A8",
  5795 => x"F800",
  5796 => x"A8A8",
  5797 => x"A8A8",
  5798 => x"A8F8",
  5799 => x"0800",
  5800 => x"C040",
  5801 => x"4070",
  5802 => x"4848",
  5803 => x"7000",
  5804 => x"8888",
  5805 => x"88E8",
  5806 => x"9898",
  5807 => x"E800",
  5808 => x"8080",
  5809 => x"80F0",
  5810 => x"8888",
  5811 => x"F000",
  5812 => x"7088",
  5813 => x"0878",
  5814 => x"0888",
  5815 => x"7000",
  5816 => x"90A8",
  5817 => x"A8E8",
  5818 => x"A8A8",
  5819 => x"9000",
  5820 => x"7888",
  5821 => x"8878",
  5822 => x"4888",
  5823 => x"8800",
  5824 => x"0000",
  5825 => x"0000",
  5826 => x"0000",
  5827 => x"0000",
  5828 => x"0000",
  5829 => x"0000",
  5830 => x"0000",
  5831 => x"0000",
  5832 => x"0000",
  5833 => x"0000",
  5834 => x"0000",
  5835 => x"0000",
  5836 => x"0000",
  5837 => x"0000",
  5838 => x"0000",
  5839 => x"0000",
  5840 => x"760F",
  5841 => x"080F",
  5842 => x"6300",
  5843 => x"6101",
  5844 => x"6002",
  5845 => x"6A03",
  5846 => x"1D00",
  5847 => x"1C01",
  5848 => x"0102",
  5849 => x"2303",
  5850 => x"0000",
  5851 => x"7500",
  5852 => x"6B01",
  5853 => x"7202",
  5854 => x"7403",
  5855 => x"0000",
  5856 => x"CFF1",
  5857 => x"300E",
  5858 => x"C7C1",
  5859 => x"2832",
  5860 => x"C301",
  5861 => x"24C2",
  5862 => x"C003",
  5863 => x"2304",
  5864 => x"C007",
  5865 => x"2008",
  5866 => x"C00F",
  5867 => x"2010",
  5868 => x"801F",
  5869 => x"4020",
  5870 => x"803F",
  5871 => x"4040",
  5872 => x"807F",
  5873 => x"4080",
  5874 => x"80FF",
  5875 => x"4100",
  5876 => x"81FF",
  5877 => x"4200",
  5878 => x"03FF",
  5879 => x"8400",
  5880 => x"07FF",
  5881 => x"8800",
  5882 => x"0FFF",
  5883 => x"9000",
  5884 => x"1FFF",
  5885 => x"A000",
  5886 => x"3FFF",
  5887 => x"C000",
  5888 => x"E3F1",
  5889 => x"1C0E",
  5890 => x"E1C1",
  5891 => x"1232",
  5892 => x"E083",
  5893 => x"1144",
  5894 => x"E003",
  5895 => x"1084",
  5896 => x"E007",
  5897 => x"1008",
  5898 => x"F007",
  5899 => x"0808",
  5900 => x"F00F",
  5901 => x"0810",
  5902 => x"F00F",
  5903 => x"0810",
  5904 => x"F01F",
  5905 => x"0820",
  5906 => x"F01F",
  5907 => x"0820",
  5908 => x"F03F",
  5909 => x"0840",
  5910 => x"F83F",
  5911 => x"0440",
  5912 => x"F87F",
  5913 => x"0480",
  5914 => x"F87F",
  5915 => x"0480",
  5916 => x"F8FF",
  5917 => x"0500",
  5918 => x"F9FF",
  5919 => x"0600",
  5920 => x"8FF1",
  5921 => x"700E",
  5922 => x"83C1",
  5923 => x"4C32",
  5924 => x"8181",
  5925 => x"4242",
  5926 => x"8001",
  5927 => x"4182",
  5928 => x"8001",
  5929 => x"4002",
  5930 => x"C003",
  5931 => x"2004",
  5932 => x"C003",
  5933 => x"2004",
  5934 => x"C003",
  5935 => x"2004",
  5936 => x"E007",
  5937 => x"1008",
  5938 => x"E007",
  5939 => x"1008",
  5940 => x"F00F",
  5941 => x"0810",
  5942 => x"F00F",
  5943 => x"0810",
  5944 => x"F81F",
  5945 => x"0420",
  5946 => x"F81F",
  5947 => x"0420",
  5948 => x"FC3F",
  5949 => x"0240",
  5950 => x"FE7F",
  5951 => x"0180",
  5952 => x"8FC7",
  5953 => x"7038",
  5954 => x"8387",
  5955 => x"4C48",
  5956 => x"C107",
  5957 => x"2288",
  5958 => x"C007",
  5959 => x"2108",
  5960 => x"E007",
  5961 => x"1008",
  5962 => x"E00F",
  5963 => x"1010",
  5964 => x"F00F",
  5965 => x"0810",
  5966 => x"F00F",
  5967 => x"0810",
  5968 => x"F80F",
  5969 => x"0410",
  5970 => x"F80F",
  5971 => x"0410",
  5972 => x"FC0F",
  5973 => x"0210",
  5974 => x"FC1F",
  5975 => x"0220",
  5976 => x"FE1F",
  5977 => x"0120",
  5978 => x"FE1F",
  5979 => x"0120",
  5980 => x"FF1F",
  5981 => x"00A0",
  5982 => x"FF9F",
  5983 => x"0060",
  5984 => x"8FF3",
  5985 => x"700C",
  5986 => x"83E3",
  5987 => x"4C14",
  5988 => x"80C3",
  5989 => x"4324",
  5990 => x"C003",
  5991 => x"20C4",
  5992 => x"E003",
  5993 => x"1004",
  5994 => x"F003",
  5995 => x"0804",
  5996 => x"F801",
  5997 => x"0402",
  5998 => x"FC01",
  5999 => x"0202",
  6000 => x"FE01",
  6001 => x"0102",
  6002 => x"FF01",
  6003 => x"0082",
  6004 => x"FF81",
  6005 => x"0042",
  6006 => x"FFC0",
  6007 => x"0021",
  6008 => x"FFE0",
  6009 => x"0011",
  6010 => x"FFF0",
  6011 => x"0009",
  6012 => x"FFF8",
  6013 => x"0005",
  6014 => x"FFFC",
  6015 => x"0003",
  6016 => x"180C",
  6017 => x"06FF",
  6018 => x"060C",
  6019 => x"1800",
  6020 => x"1038",
  6021 => x"7CD6",
  6022 => x"9210",
  6023 => x"1010",
  6024 => x"1010",
  6025 => x"1092",
  6026 => x"D67C",
  6027 => x"3810",
  6028 => x"0000",
  6029 => x"0000",
  6030 => x"0000",
  6031 => x"0000",
  6032 => x"00FC",
  6033 => x"FEFF",
  6034 => x"FFFE",
  6035 => x"FC00",
  6036 => x"003F",
  6037 => x"7FFF",
  6038 => x"FF7F",
  6039 => x"3F00",
  6040 => x"00FF",
  6041 => x"FFFF",
  6042 => x"FFFF",
  6043 => x"FF00",
  6044 => x"0000",
  6045 => x"0000",
  6046 => x"0000",
  6047 => x"0000",
  6048 => x"0000",
  6049 => x"0000",
  6050 => x"0000",
  6051 => x"0000",
  6052 => x"5061",
  6053 => x"7065",
  6054 => x"7250",
  6055 => x"6C61",
  6056 => x"6E65",
  6057 => x"0000",
  6058 => x"6D2F",
  6059 => x"7300",
  6060 => x"0000",
  6061 => x"0000",
  6062 => x"0000",
  6063 => x"0000",
  6064 => x"0000",
  6065 => x"0000",
  6066 => x"0000",
  6067 => x"0000",
  6068 => x"0000",
  6069 => x"0000",
  6070 => x"0000",
  6071 => x"0000",
  6072 => x"0000",
  6073 => x"0000",
  6074 => x"0000",
  6075 => x"0000",
  6076 => x"0000",
  6077 => x"0000",
  6078 => x"0000",
  6079 => x"0000",
  6080 => x"0000",
  6081 => x"0000",
  6082 => x"0000",
  6083 => x"0000",
  6084 => x"0000",
  6085 => x"0000",
  6086 => x"0000",
  6087 => x"0000",
  6088 => x"0000",
  6089 => x"0000",
  6090 => x"0000",
  6091 => x"0000",
  6092 => x"0000",
  6093 => x"0000",
  6094 => x"0000",
  6095 => x"0000",
  6096 => x"0000",
  6097 => x"0000",
  6098 => x"0000",
  6099 => x"0000",
  6100 => x"0000",
  6101 => x"0000",
  6102 => x"0000",
  6103 => x"0000",
  6104 => x"0000",
  6105 => x"0000",
  6106 => x"0000",
  6107 => x"0000",
  6108 => x"0000",
  6109 => x"0000",
  6110 => x"0000",
  6111 => x"0000",
  6112 => x"0000",
  6113 => x"0000",
  6114 => x"0000",
  6115 => x"0000",
  6116 => x"0000",
  6117 => x"0000",
  6118 => x"0000",
  6119 => x"0000",
  6120 => x"0000",
  6121 => x"0000",
  6122 => x"0000",
  6123 => x"0000",
  6124 => x"0000",
  6125 => x"0000",
  6126 => x"0000",
  6127 => x"0000",
  6128 => x"0000",
  6129 => x"0000",
  6130 => x"0000",
  6131 => x"0000",
  6132 => x"0000",
  6133 => x"0000",
  6134 => x"0000",
  6135 => x"0000",
  6136 => x"0000",
  6137 => x"0000",
  6138 => x"0000",
  6139 => x"0000",
  6140 => x"0000",
  6141 => x"0000",
  6142 => x"0000",
  6143 => x"0000",
  6144 => x"0000",
  6145 => x"0000",
  6146 => x"0000",
  6147 => x"0000",
  6148 => x"0000",
  6149 => x"0000",
  6150 => x"0000",
  6151 => x"0000",
  6152 => x"0000",
  6153 => x"0000",
  6154 => x"0000",
  6155 => x"0000",
  6156 => x"0000",
  6157 => x"0000",
  6158 => x"0000",
  6159 => x"0000",
  6160 => x"0000",
  6161 => x"0000",
  6162 => x"0000",
  6163 => x"0000",
  6164 => x"0000",
  6165 => x"0000",
  6166 => x"0000",
  6167 => x"0000",
  6168 => x"0000",
  6169 => x"0000",
  6170 => x"0000",
  6171 => x"0000",
  6172 => x"0000",
  6173 => x"0000",
  6174 => x"0000",
  6175 => x"0000",
  6176 => x"0000",
  6177 => x"0000",
  6178 => x"0000",
  6179 => x"0000",
  6180 => x"0000",
  6181 => x"0000",
  6182 => x"0000",
  6183 => x"0000",
  6184 => x"0000",
  6185 => x"0000",
  6186 => x"0000",
  6187 => x"0000",
  6188 => x"0000",
  6189 => x"0000",
  6190 => x"0000",
  6191 => x"0000",
  6192 => x"0000",
  6193 => x"0000",
  6194 => x"0000",
  6195 => x"0000",
  6196 => x"0000",
  6197 => x"0000",
  6198 => x"0000",
  6199 => x"0000",
  6200 => x"0000",
  6201 => x"0000",
  6202 => x"0000",
  6203 => x"0000",
  6204 => x"0000",
  6205 => x"0000",
  6206 => x"0000",
  6207 => x"0000",
  6208 => x"0000",
  6209 => x"0000",
  6210 => x"0000",
  6211 => x"0000",
  6212 => x"0000",
  6213 => x"0000",
  6214 => x"0000",
  6215 => x"0000",
  6216 => x"0000",
  6217 => x"0000",
  6218 => x"0000",
  6219 => x"0000",
  6220 => x"0000",
  6221 => x"0000",
  6222 => x"0000",
  6223 => x"0000",
  6224 => x"0000",
  6225 => x"0000",
  6226 => x"0000",
  6227 => x"0000",
  6228 => x"0000",
  6229 => x"0000",
  6230 => x"0000",
  6231 => x"0000",
  6232 => x"0000",
  6233 => x"0000",
  6234 => x"0000",
  6235 => x"0000",
  6236 => x"0000",
  6237 => x"0000",
  6238 => x"0000",
  6239 => x"0000",
  6240 => x"0000",
  6241 => x"0000",
  6242 => x"0000",
  6243 => x"0000",
  6244 => x"0000",
  6245 => x"0000",
  6246 => x"0000",
  6247 => x"0000",
  6248 => x"0000",
  6249 => x"0000",
  6250 => x"0000",
  6251 => x"0000",
  6252 => x"0000",
  6253 => x"0000",
  6254 => x"0000",
  6255 => x"0000",
  6256 => x"0000",
  6257 => x"0000",
  6258 => x"0000",
  6259 => x"0000",
  6260 => x"0000",
  6261 => x"0000",
  6262 => x"0000",
  6263 => x"0000",
  6264 => x"0000",
  6265 => x"0000",
  6266 => x"0000",
  6267 => x"0000",
  6268 => x"0000",
  6269 => x"0000",
  6270 => x"0000",
  6271 => x"0000",
  6272 => x"0000",
  6273 => x"0000",
  6274 => x"0000",
  6275 => x"0000",
  6276 => x"0000",
  6277 => x"0000",
  6278 => x"0000",
  6279 => x"0000",
  6280 => x"0000",
  6281 => x"0000",
  6282 => x"0000",
  6283 => x"0000",
  6284 => x"0000",
  6285 => x"0000",
  6286 => x"0000",
  6287 => x"0000",
  6288 => x"0000",
  6289 => x"0000",
  6290 => x"0000",
  6291 => x"0000",
  6292 => x"0000",
  6293 => x"0000",
  6294 => x"0000",
  6295 => x"0000",
  6296 => x"0000",
  6297 => x"0000",
  6298 => x"0000",
  6299 => x"0000",
  6300 => x"0000",
  6301 => x"0000",
  6302 => x"0000",
  6303 => x"0000",
  6304 => x"0000",
  6305 => x"0000",
  6306 => x"0000",
  6307 => x"0000",
  6308 => x"0000",
  6309 => x"0000",
  6310 => x"0000",
  6311 => x"0000",
  6312 => x"0000",
  6313 => x"0000",
  6314 => x"0000",
  6315 => x"0000",
  6316 => x"0000",
  6317 => x"0000",
  6318 => x"0000",
  6319 => x"0000",
  6320 => x"0000",
  6321 => x"0000",
  6322 => x"0000",
  6323 => x"0000",
  6324 => x"0000",
  6325 => x"0000",
  6326 => x"0000",
  6327 => x"0000",
  6328 => x"0000",
  6329 => x"0000",
  6330 => x"0000",
  6331 => x"0000",
  6332 => x"0000",
  6333 => x"0000",
  6334 => x"0000",
  6335 => x"0000",
  6336 => x"0000",
  6337 => x"0000",
  6338 => x"0000",
  6339 => x"0000",
  6340 => x"0000",
  6341 => x"0000",
  6342 => x"0000",
  6343 => x"0000",
  6344 => x"0000",
  6345 => x"0000",
  6346 => x"0000",
  6347 => x"0000",
  6348 => x"0000",
  6349 => x"0000",
  6350 => x"0000",
  6351 => x"0000",
  6352 => x"0000",
  6353 => x"0000",
  6354 => x"0000",
  6355 => x"0000",
  6356 => x"0000",
  6357 => x"0000",
  6358 => x"0000",
  6359 => x"0000",
  6360 => x"0000",
  6361 => x"0000",
  6362 => x"0000",
  6363 => x"0000",
  6364 => x"0000",
  6365 => x"0000",
  6366 => x"0000",
  6367 => x"0000",
  6368 => x"0000",
  6369 => x"0000",
  6370 => x"0000",
  6371 => x"0000",
  6372 => x"0000",
  6373 => x"0000",
  6374 => x"0000",
  6375 => x"0000",
  6376 => x"0000",
  6377 => x"0000",
  6378 => x"0000",
  6379 => x"0000",
  6380 => x"0000",
  6381 => x"0000",
  6382 => x"0000",
  6383 => x"0000",
  6384 => x"0000",
  6385 => x"0000",
  6386 => x"0000",
  6387 => x"0000",
  6388 => x"0000",
  6389 => x"0000",
  6390 => x"0000",
  6391 => x"0000",
  6392 => x"0000",
  6393 => x"0000",
  6394 => x"0000",
  6395 => x"0000",
  6396 => x"0000",
  6397 => x"0000",
  6398 => x"0000",
  6399 => x"0000",
  6400 => x"0000",
  6401 => x"0000",
  6402 => x"0000",
  6403 => x"0000",
  6404 => x"0000",
  6405 => x"0000",
  6406 => x"0000",
  6407 => x"0000",
  6408 => x"0000",
  6409 => x"0000",
  6410 => x"0000",
  6411 => x"0000",
  6412 => x"0000",
  6413 => x"0000",
  6414 => x"0000",
  6415 => x"0000",
  6416 => x"0000",
  6417 => x"0000",
  6418 => x"0000",
  6419 => x"0000",
  6420 => x"0000",
  6421 => x"0000",
  6422 => x"0000",
  6423 => x"0000",
  6424 => x"0000",
  6425 => x"0000",
  6426 => x"0000",
  6427 => x"0000",
  6428 => x"0000",
  6429 => x"0000",
  6430 => x"0000",
  6431 => x"0000",
  6432 => x"0000",
  6433 => x"0000",
  6434 => x"0000",
  6435 => x"0000",
  6436 => x"0000",
  6437 => x"0000",
  6438 => x"0000",
  6439 => x"0000",
  6440 => x"0000",
  6441 => x"0000",
  6442 => x"0000",
  6443 => x"0000",
  6444 => x"0000",
  6445 => x"0000",
  6446 => x"0000",
  6447 => x"0000",
  6448 => x"0000",
  6449 => x"0000",
  6450 => x"0000",
  6451 => x"0000",
  6452 => x"0000",
  6453 => x"0000",
  6454 => x"0000",
  6455 => x"0000",
  6456 => x"0000",
  6457 => x"0000",
  6458 => x"0000",
  6459 => x"0000",
  6460 => x"0000",
  6461 => x"0000",
  6462 => x"0000",
  6463 => x"0000",
  6464 => x"0000",
  6465 => x"0000",
  6466 => x"0000",
  6467 => x"0000",
  6468 => x"0000",
  6469 => x"0000",
  6470 => x"0000",
  6471 => x"0000",
  6472 => x"0000",
  6473 => x"0000",
  6474 => x"0000",
  6475 => x"0000",
  6476 => x"0000",
  6477 => x"0000",
  6478 => x"0000",
  6479 => x"0000",
  6480 => x"0000",
  6481 => x"0000",
  6482 => x"0000",
  6483 => x"0000",
  6484 => x"0000",
  6485 => x"0000",
  6486 => x"0000",
  6487 => x"0000",
  6488 => x"0000",
  6489 => x"0000",
  6490 => x"0000",
  6491 => x"0000",
  6492 => x"0000",
  6493 => x"0000",
  6494 => x"0000",
  6495 => x"0000",
  6496 => x"0000",
  6497 => x"0000",
  6498 => x"0000",
  6499 => x"0000",
  6500 => x"0000",
  6501 => x"0000",
  6502 => x"0000",
  6503 => x"0000",
  6504 => x"0000",
  6505 => x"0000",
  6506 => x"0000",
  6507 => x"0000",
  6508 => x"0000",
  6509 => x"0000",
  6510 => x"0000",
  6511 => x"0000",
  6512 => x"0000",
  6513 => x"0000",
  6514 => x"0000",
  6515 => x"0000",
  6516 => x"0000",
  6517 => x"0000",
  6518 => x"0000",
  6519 => x"0000",
  6520 => x"0000",
  6521 => x"0000",
  6522 => x"0000",
  6523 => x"0000",
  6524 => x"0000",
  6525 => x"0000",
  6526 => x"0000",
  6527 => x"0000",
  6528 => x"0000",
  6529 => x"0000",
  6530 => x"0000",
  6531 => x"0000",
  6532 => x"0000",
  6533 => x"0000",
  6534 => x"0000",
  6535 => x"0000",
  6536 => x"0000",
  6537 => x"0000",
  6538 => x"0000",
  6539 => x"0000",
  6540 => x"0000",
  6541 => x"0000",
  6542 => x"0000",
  6543 => x"0000",
  6544 => x"0000",
  6545 => x"0000",
  6546 => x"0000",
  6547 => x"0000",
  6548 => x"0000",
  6549 => x"0000",
  6550 => x"0000",
  6551 => x"0000",
  6552 => x"0000",
  6553 => x"0000",
  6554 => x"0000",
  6555 => x"0000",
  6556 => x"0000",
  6557 => x"0000",
  6558 => x"0000",
  6559 => x"0000",
  6560 => x"0000",
  6561 => x"0000",
  6562 => x"0000",
  6563 => x"0000",
  6564 => x"0000",
  6565 => x"0000",
  6566 => x"0000",
  6567 => x"0000",
  6568 => x"0000",
  6569 => x"0000",
  6570 => x"0000",
  6571 => x"0000",
  6572 => x"0000",
  6573 => x"0000",
  6574 => x"0000",
  6575 => x"0000",
  6576 => x"0000",
  6577 => x"0000",
  6578 => x"0000",
  6579 => x"0000",
  6580 => x"0000",
  6581 => x"0000",
  6582 => x"0000",
  6583 => x"0000",
  6584 => x"0000",
  6585 => x"0000",
  6586 => x"0000",
  6587 => x"0000",
  6588 => x"0000",
  6589 => x"0000",
  6590 => x"0000",
  6591 => x"0000",
  6592 => x"0000",
  6593 => x"0000",
  6594 => x"0000",
  6595 => x"0000",
  6596 => x"0000",
  6597 => x"0000",
  6598 => x"0000",
  6599 => x"0000",
  6600 => x"0000",
  6601 => x"0000",
  6602 => x"0000",
  6603 => x"0000",
  6604 => x"0000",
  6605 => x"0000",
  6606 => x"0000",
  6607 => x"0000",
  6608 => x"0000",
  6609 => x"0000",
  6610 => x"0000",
  6611 => x"0000",
  6612 => x"0000",
  6613 => x"0000",
  6614 => x"0000",
  6615 => x"0000",
  6616 => x"0000",
  6617 => x"0000",
  6618 => x"0000",
  6619 => x"0000",
  6620 => x"0000",
  6621 => x"0000",
  6622 => x"0000",
  6623 => x"0000",
  6624 => x"0000",
  6625 => x"0000",
  6626 => x"0000",
  6627 => x"0000",
  6628 => x"0000",
  6629 => x"0000",
  6630 => x"0000",
  6631 => x"0000",
  6632 => x"0000",
  6633 => x"0000",
  6634 => x"0000",
  6635 => x"0000",
  6636 => x"0000",
  6637 => x"0000",
  6638 => x"0000",
  6639 => x"0000",
  6640 => x"0000",
  6641 => x"0000",
  6642 => x"0000",
  6643 => x"0000",
  6644 => x"0000",
  6645 => x"0000",
  6646 => x"0000",
  6647 => x"0000",
  6648 => x"0000",
  6649 => x"0000",
  6650 => x"0000",
  6651 => x"0000",
  6652 => x"0000",
  6653 => x"0000",
  6654 => x"0000",
  6655 => x"0000",
  6656 => x"0000",
  6657 => x"0000",
  6658 => x"0000",
  6659 => x"0000",
  6660 => x"0000",
  6661 => x"0000",
  6662 => x"0000",
  6663 => x"0000",
  6664 => x"0000",
  6665 => x"0000",
  6666 => x"0000",
  6667 => x"0000",
  6668 => x"0000",
  6669 => x"0000",
  6670 => x"0000",
  6671 => x"0000",
  6672 => x"0000",
  6673 => x"0000",
  6674 => x"0000",
  6675 => x"0000",
  6676 => x"0000",
  6677 => x"0000",
  6678 => x"0000",
  6679 => x"0000",
  6680 => x"0000",
  6681 => x"0000",
  6682 => x"0000",
  6683 => x"0000",
  6684 => x"0000",
  6685 => x"0000",
  6686 => x"0000",
  6687 => x"0000",
  6688 => x"0000",
  6689 => x"0000",
  6690 => x"0000",
  6691 => x"0000",
  6692 => x"0000",
  6693 => x"0000",
  6694 => x"0000",
  6695 => x"0000",
  6696 => x"0000",
  6697 => x"0000",
  6698 => x"0000",
  6699 => x"0000",
  6700 => x"0000",
  6701 => x"0000",
  6702 => x"0000",
  6703 => x"0000",
  6704 => x"0000",
  6705 => x"0000",
  6706 => x"0000",
  6707 => x"0000",
  6708 => x"0000",
  6709 => x"0000",
  6710 => x"0000",
  6711 => x"0000",
  6712 => x"0000",
  6713 => x"0000",
  6714 => x"0000",
  6715 => x"0000",
  6716 => x"0000",
  6717 => x"0000",
  6718 => x"0000",
  6719 => x"0000",
  6720 => x"0000",
  6721 => x"0000",
  6722 => x"0000",
  6723 => x"0000",
  6724 => x"0000",
  6725 => x"0000",
  6726 => x"0000",
  6727 => x"0000",
  6728 => x"0000",
  6729 => x"0000",
  6730 => x"0000",
  6731 => x"0000",
  6732 => x"0000",
  6733 => x"0000",
  6734 => x"0000",
  6735 => x"0000",
  6736 => x"0000",
  6737 => x"0000",
  6738 => x"0000",
  6739 => x"0000",
  6740 => x"0000",
  6741 => x"0000",
  6742 => x"0000",
  6743 => x"0000",
  6744 => x"0000",
  6745 => x"0000",
  6746 => x"0000",
  6747 => x"0000",
  6748 => x"0000",
  6749 => x"0000",
  6750 => x"0000",
  6751 => x"0000",
  6752 => x"0000",
  6753 => x"0000",
  6754 => x"0000",
  6755 => x"0000",
  6756 => x"0000",
  6757 => x"0000",
  6758 => x"0000",
  6759 => x"0000",
  6760 => x"0000",
  6761 => x"0000",
  6762 => x"0000",
  6763 => x"0000",
  6764 => x"0000",
  6765 => x"0000",
  6766 => x"0000",
  6767 => x"0000",
  6768 => x"0000",
  6769 => x"0000",
  6770 => x"0000",
  6771 => x"0000",
  6772 => x"0000",
  6773 => x"0000",
  6774 => x"0000",
  6775 => x"0000",
  6776 => x"0000",
  6777 => x"0000",
  6778 => x"0000",
  6779 => x"0000",
  6780 => x"0000",
  6781 => x"0000",
  6782 => x"0000",
  6783 => x"0000",
  6784 => x"0000",
  6785 => x"0000",
  6786 => x"0000",
  6787 => x"0000",
  6788 => x"0000",
  6789 => x"0000",
  6790 => x"0000",
  6791 => x"0000",
  6792 => x"0000",
  6793 => x"0000",
  6794 => x"0000",
  6795 => x"0000",
  6796 => x"0000",
  6797 => x"0000",
  6798 => x"0000",
  6799 => x"0000",
  6800 => x"0000",
  6801 => x"0000",
  6802 => x"0000",
  6803 => x"0000",
  6804 => x"0000",
  6805 => x"0000",
  6806 => x"0000",
  6807 => x"0000",
  6808 => x"0000",
  6809 => x"0000",
  6810 => x"0000",
  6811 => x"0000",
  6812 => x"0000",
  6813 => x"0000",
  6814 => x"0000",
  6815 => x"0000",
  6816 => x"0000",
  6817 => x"0000",
  6818 => x"0000",
  6819 => x"0000",
  6820 => x"0000",
  6821 => x"0000",
  6822 => x"0000",
  6823 => x"0000",
  6824 => x"0000",
  6825 => x"0000",
  6826 => x"0000",
  6827 => x"0000",
  6828 => x"0000",
  6829 => x"0000",
  6830 => x"0000",
  6831 => x"0000",
  6832 => x"0000",
  6833 => x"0000",
  6834 => x"0000",
  6835 => x"0000",
  6836 => x"0000",
  6837 => x"0000",
  6838 => x"0000",
  6839 => x"0000",
  6840 => x"0000",
  6841 => x"0000",
  6842 => x"0000",
  6843 => x"0000",
  6844 => x"0000",
  6845 => x"0000",
  6846 => x"0000",
  6847 => x"0000",
  6848 => x"0000",
  6849 => x"0000",
  6850 => x"0000",
  6851 => x"0000",
  6852 => x"0000",
  6853 => x"0000",
  6854 => x"0000",
  6855 => x"0000",
  6856 => x"0000",
  6857 => x"0000",
  6858 => x"0000",
  6859 => x"0000",
  6860 => x"0000",
  6861 => x"0000",
  6862 => x"0000",
  6863 => x"0000",
  6864 => x"0000",
  6865 => x"0000",
  6866 => x"0000",
  6867 => x"0000",
  6868 => x"0000",
  6869 => x"0000",
  6870 => x"0000",
  6871 => x"0000",
  6872 => x"0000",
  6873 => x"0000",
  6874 => x"0000",
  6875 => x"0000",
  6876 => x"0000",
  6877 => x"0000",
  6878 => x"0000",
  6879 => x"0000",
  6880 => x"0000",
  6881 => x"0000",
  6882 => x"0000",
  6883 => x"0000",
  6884 => x"0000",
  6885 => x"0000",
  6886 => x"0000",
  6887 => x"0000",
  6888 => x"0000",
  6889 => x"0000",
  6890 => x"0000",
  6891 => x"0000",
  6892 => x"0000",
  6893 => x"0000",
  6894 => x"0000",
  6895 => x"0000",
  6896 => x"0000",
  6897 => x"0000",
  6898 => x"0000",
  6899 => x"0000",
  6900 => x"0000",
  6901 => x"0000",
  6902 => x"0000",
  6903 => x"0000",
  6904 => x"0000",
  6905 => x"0000",
  6906 => x"0000",
  6907 => x"0000",
  6908 => x"0000",
  6909 => x"0000",
  6910 => x"0000",
  6911 => x"0000",
  6912 => x"0000",
  6913 => x"0000",
  6914 => x"0000",
  6915 => x"0000",
  6916 => x"0000",
  6917 => x"0000",
  6918 => x"0000",
  6919 => x"0000",
  6920 => x"0000",
  6921 => x"0000",
  6922 => x"0000",
  6923 => x"0000",
  6924 => x"0000",
  6925 => x"0000",
  6926 => x"0000",
  6927 => x"0000",
  6928 => x"0000",
  6929 => x"0000",
  6930 => x"0000",
  6931 => x"0000",
  6932 => x"0000",
  6933 => x"0000",
  6934 => x"0000",
  6935 => x"0000",
  6936 => x"0000",
  6937 => x"0000",
  6938 => x"0000",
  6939 => x"0000",
  6940 => x"0000",
  6941 => x"0000",
  6942 => x"0000",
  6943 => x"0000",
  6944 => x"0000",
  6945 => x"0000",
  6946 => x"0000",
  6947 => x"0000",
  6948 => x"0000",
  6949 => x"0000",
  6950 => x"0000",
  6951 => x"0000",
  6952 => x"0000",
  6953 => x"0000",
  6954 => x"0000",
  6955 => x"0000",
  6956 => x"0000",
  6957 => x"0000",
  6958 => x"0000",
  6959 => x"0000",
  6960 => x"0000",
  6961 => x"0000",
  6962 => x"0000",
  6963 => x"0000",
  6964 => x"0000",
  6965 => x"0000",
  6966 => x"0000",
  6967 => x"0000",
  6968 => x"0000",
  6969 => x"0000",
  6970 => x"0000",
  6971 => x"0000",
  6972 => x"0000",
  6973 => x"0000",
  6974 => x"0000",
  6975 => x"0000",
  6976 => x"0000",
  6977 => x"0000",
  6978 => x"0000",
  6979 => x"0000",
  6980 => x"0000",
  6981 => x"0000",
  6982 => x"0000",
  6983 => x"0000",
  6984 => x"0000",
  6985 => x"0000",
  6986 => x"0000",
  6987 => x"0000",
  6988 => x"0000",
  6989 => x"0000",
  6990 => x"0000",
  6991 => x"0000",
  6992 => x"0000",
  6993 => x"0000",
  6994 => x"0000",
  6995 => x"0000",
  6996 => x"0000",
  6997 => x"0000",
  6998 => x"0000",
  6999 => x"0000",
  7000 => x"0000",
  7001 => x"0000",
  7002 => x"0000",
  7003 => x"0000",
  7004 => x"0000",
  7005 => x"0000",
  7006 => x"0000",
  7007 => x"0000",
  7008 => x"0000",
  7009 => x"0000",
  7010 => x"0000",
  7011 => x"0000",
  7012 => x"0000",
  7013 => x"0000",
  7014 => x"0000",
  7015 => x"0000",
  7016 => x"0000",
  7017 => x"0000",
  7018 => x"0000",
  7019 => x"0000",
  7020 => x"0000",
  7021 => x"0000",
  7022 => x"0000",
  7023 => x"0000",
  7024 => x"0000",
  7025 => x"0000",
  7026 => x"0000",
  7027 => x"0000",
  7028 => x"0000",
  7029 => x"0000",
  7030 => x"0000",
  7031 => x"0000",
  7032 => x"0000",
  7033 => x"0000",
  7034 => x"0000",
  7035 => x"0000",
  7036 => x"0000",
  7037 => x"0000",
  7038 => x"0000",
  7039 => x"0000",
  7040 => x"0000",
  7041 => x"0000",
  7042 => x"0000",
  7043 => x"0000",
  7044 => x"0000",
  7045 => x"0000",
  7046 => x"0000",
  7047 => x"0000",
  7048 => x"0000",
  7049 => x"0000",
  7050 => x"0000",
  7051 => x"0000",
  7052 => x"0000",
  7053 => x"0000",
  7054 => x"0000",
  7055 => x"0000",
  7056 => x"0000",
  7057 => x"0000",
  7058 => x"0000",
  7059 => x"0000",
  7060 => x"0000",
  7061 => x"0000",
  7062 => x"0000",
  7063 => x"0000",
  7064 => x"0000",
  7065 => x"0000",
  7066 => x"0000",
  7067 => x"0000",
  7068 => x"0000",
  7069 => x"0000",
  7070 => x"0000",
  7071 => x"0000",
  7072 => x"0000",
  7073 => x"0000",
  7074 => x"0000",
  7075 => x"0000",
  7076 => x"0000",
  7077 => x"0000",
  7078 => x"0000",
  7079 => x"0000",
  7080 => x"0000",
  7081 => x"0000",
  7082 => x"0000",
  7083 => x"0000",
  7084 => x"0000",
  7085 => x"0000",
  7086 => x"0000",
  7087 => x"0000",
  7088 => x"0000",
  7089 => x"0000",
  7090 => x"0000",
  7091 => x"0000",
  7092 => x"0000",
  7093 => x"0000",
  7094 => x"0000",
  7095 => x"0000",
  7096 => x"0000",
  7097 => x"0000",
  7098 => x"0000",
  7099 => x"0000",
  7100 => x"0000",
  7101 => x"0000",
  7102 => x"0000",
  7103 => x"0000",
  7104 => x"0000",
  7105 => x"0000",
  7106 => x"0000",
  7107 => x"0000",
  7108 => x"0000",
  7109 => x"0000",
  7110 => x"0000",
  7111 => x"0000",
  7112 => x"0000",
  7113 => x"0000",
  7114 => x"0000",
  7115 => x"0000",
  7116 => x"0000",
  7117 => x"0000",
  7118 => x"0000",
  7119 => x"0000",
  7120 => x"0000",
  7121 => x"0000",
  7122 => x"0000",
  7123 => x"0000",
  7124 => x"0000",
  7125 => x"0000",
  7126 => x"0000",
  7127 => x"0000",
  7128 => x"0000",
  7129 => x"0000",
  7130 => x"0000",
  7131 => x"0000",
  7132 => x"0000",
  7133 => x"0000",
  7134 => x"0000",
  7135 => x"0000",
  7136 => x"0000",
  7137 => x"0000",
  7138 => x"0000",
  7139 => x"0000",
  7140 => x"0000",
  7141 => x"0000",
  7142 => x"0000",
  7143 => x"0000",
  7144 => x"0000",
  7145 => x"0000",
  7146 => x"0000",
  7147 => x"0000",
  7148 => x"0000",
  7149 => x"0000",
  7150 => x"0000",
  7151 => x"0000",
  7152 => x"0000",
  7153 => x"0000",
  7154 => x"0000",
  7155 => x"0000",
  7156 => x"0000",
  7157 => x"0000",
  7158 => x"0000",
  7159 => x"0000",
  7160 => x"0000",
  7161 => x"0000",
  7162 => x"0000",
  7163 => x"0000",
  7164 => x"0000",
  7165 => x"0000",
  7166 => x"0000",
  7167 => x"0000",
  7168 => x"0000",
  7169 => x"0000",
  7170 => x"0000",
  7171 => x"0000",
  7172 => x"0000",
  7173 => x"0000",
  7174 => x"0000",
  7175 => x"0000",
  7176 => x"0000",
  7177 => x"0000",
  7178 => x"0000",
  7179 => x"0000",
  7180 => x"0000",
  7181 => x"0000",
  7182 => x"0000",
  7183 => x"0000",
  7184 => x"0000",
  7185 => x"0000",
  7186 => x"0000",
  7187 => x"0000",
  7188 => x"0000",
  7189 => x"0000",
  7190 => x"0000",
  7191 => x"0000",
  7192 => x"0000",
  7193 => x"0000",
  7194 => x"0000",
  7195 => x"0000",
  7196 => x"0000",
  7197 => x"0000",
  7198 => x"0000",
  7199 => x"0000",
  7200 => x"0000",
  7201 => x"0000",
  7202 => x"0000",
  7203 => x"0000",
  7204 => x"0000",
  7205 => x"0000",
  7206 => x"0000",
  7207 => x"0000",
  7208 => x"0000",
  7209 => x"0000",
  7210 => x"0000",
  7211 => x"0000",
  7212 => x"0000",
  7213 => x"0000",
  7214 => x"0000",
  7215 => x"0000",
  7216 => x"0000",
  7217 => x"0000",
  7218 => x"0000",
  7219 => x"0000",
  7220 => x"0000",
  7221 => x"0000",
  7222 => x"0000",
  7223 => x"0000",
  7224 => x"0000",
  7225 => x"0000",
  7226 => x"0000",
  7227 => x"0000",
  7228 => x"0000",
  7229 => x"0000",
  7230 => x"0000",
  7231 => x"0000",
  7232 => x"0000",
  7233 => x"0000",
  7234 => x"0000",
  7235 => x"0000",
  7236 => x"0000",
  7237 => x"0000",
  7238 => x"0000",
  7239 => x"0000",
  7240 => x"0000",
  7241 => x"0000",
  7242 => x"0000",
  7243 => x"0000",
  7244 => x"0000",
  7245 => x"0000",
  7246 => x"0000",
  7247 => x"0000",
  7248 => x"0000",
  7249 => x"0000",
  7250 => x"0000",
  7251 => x"0000",
  7252 => x"0000",
  7253 => x"0000",
  7254 => x"0000",
  7255 => x"0000",
  7256 => x"0000",
  7257 => x"0000",
  7258 => x"0000",
  7259 => x"0000",
  7260 => x"0000",
  7261 => x"0000",
  7262 => x"0000",
  7263 => x"0000",
  7264 => x"0000",
  7265 => x"0000",
  7266 => x"0000",
  7267 => x"0000",
  7268 => x"0000",
  7269 => x"0000",
  7270 => x"0000",
  7271 => x"0000",
  7272 => x"0000",
  7273 => x"0000",
  7274 => x"0000",
  7275 => x"0000",
  7276 => x"0000",
  7277 => x"0000",
  7278 => x"0000",
  7279 => x"0000",
  7280 => x"0000",
  7281 => x"0000",
  7282 => x"0000",
  7283 => x"0000",
  7284 => x"0000",
  7285 => x"0000",
  7286 => x"0000",
  7287 => x"0000",
  7288 => x"0000",
  7289 => x"0000",
  7290 => x"0000",
  7291 => x"0000",
  7292 => x"0000",
  7293 => x"0000",
  7294 => x"0000",
  7295 => x"0000",
  7296 => x"0000",
  7297 => x"0000",
  7298 => x"0000",
  7299 => x"0000",
  7300 => x"0000",
  7301 => x"0000",
  7302 => x"0000",
  7303 => x"0000",
  7304 => x"0000",
  7305 => x"0000",
  7306 => x"0000",
  7307 => x"0000",
  7308 => x"0000",
  7309 => x"0000",
  7310 => x"0000",
  7311 => x"0000",
  7312 => x"0000",
  7313 => x"0000",
  7314 => x"0000",
  7315 => x"0000",
  7316 => x"0000",
  7317 => x"0000",
  7318 => x"0000",
  7319 => x"0000",
  7320 => x"0000",
  7321 => x"0000",
  7322 => x"0000",
  7323 => x"0000",
  7324 => x"0000",
  7325 => x"0000",
  7326 => x"0000",
  7327 => x"0000",
  7328 => x"0000",
  7329 => x"0000",
  7330 => x"0000",
  7331 => x"0000",
  7332 => x"0000",
  7333 => x"0000",
  7334 => x"0000",
  7335 => x"0000",
  7336 => x"0000",
  7337 => x"0000",
  7338 => x"0000",
  7339 => x"0000",
  7340 => x"0000",
  7341 => x"0000",
  7342 => x"0000",
  7343 => x"0000",
  7344 => x"0000",
  7345 => x"0000",
  7346 => x"0000",
  7347 => x"0000",
  7348 => x"0000",
  7349 => x"0000",
  7350 => x"0000",
  7351 => x"0000",
  7352 => x"0000",
  7353 => x"0000",
  7354 => x"0000",
  7355 => x"0000",
  7356 => x"0000",
  7357 => x"0000",
  7358 => x"0000",
  7359 => x"0000",
  7360 => x"0000",
  7361 => x"0000",
  7362 => x"0000",
  7363 => x"0000",
  7364 => x"0000",
  7365 => x"0000",
  7366 => x"0000",
  7367 => x"0000",
  7368 => x"0000",
  7369 => x"0000",
  7370 => x"0000",
  7371 => x"0000",
  7372 => x"0000",
  7373 => x"0000",
  7374 => x"0000",
  7375 => x"0000",
  7376 => x"0000",
  7377 => x"0000",
  7378 => x"0000",
  7379 => x"0000",
  7380 => x"0000",
  7381 => x"0000",
  7382 => x"0000",
  7383 => x"0000",
  7384 => x"0000",
  7385 => x"0000",
  7386 => x"0000",
  7387 => x"0000",
  7388 => x"0000",
  7389 => x"0000",
  7390 => x"0000",
  7391 => x"0000",
  7392 => x"0000",
  7393 => x"0000",
  7394 => x"0000",
  7395 => x"0000",
  7396 => x"0000",
  7397 => x"0000",
  7398 => x"0000",
  7399 => x"0000",
  7400 => x"0000",
  7401 => x"0000",
  7402 => x"0000",
  7403 => x"0000",
  7404 => x"0000",
  7405 => x"0000",
  7406 => x"0000",
  7407 => x"0000",
  7408 => x"0000",
  7409 => x"0000",
  7410 => x"0000",
  7411 => x"0000",
  7412 => x"0000",
  7413 => x"0000",
  7414 => x"0000",
  7415 => x"0000",
  7416 => x"0000",
  7417 => x"0000",
  7418 => x"0000",
  7419 => x"0000",
  7420 => x"0000",
  7421 => x"0000",
  7422 => x"0000",
  7423 => x"0000",
  7424 => x"0000",
  7425 => x"0000",
  7426 => x"0000",
  7427 => x"0000",
  7428 => x"0000",
  7429 => x"0000",
  7430 => x"0000",
  7431 => x"0000",
  7432 => x"0000",
  7433 => x"0000",
  7434 => x"0000",
  7435 => x"0000",
  7436 => x"0000",
  7437 => x"0000",
  7438 => x"0000",
  7439 => x"0000",
  7440 => x"0000",
  7441 => x"0000",
  7442 => x"0000",
  7443 => x"0000",
  7444 => x"0000",
  7445 => x"0000",
  7446 => x"0000",
  7447 => x"0000",
  7448 => x"0000",
  7449 => x"0000",
  7450 => x"0000",
  7451 => x"0000",
  7452 => x"0000",
  7453 => x"0000",
  7454 => x"0000",
  7455 => x"0000",
  7456 => x"0000",
  7457 => x"0000",
  7458 => x"0000",
  7459 => x"0000",
  7460 => x"0000",
  7461 => x"0000",
  7462 => x"0000",
  7463 => x"0000",
  7464 => x"0000",
  7465 => x"0000",
  7466 => x"0000",
  7467 => x"0000",
  7468 => x"0000",
  7469 => x"0000",
  7470 => x"0000",
  7471 => x"0000",
  7472 => x"0000",
  7473 => x"0000",
  7474 => x"0000",
  7475 => x"0000",
  7476 => x"0000",
  7477 => x"0000",
  7478 => x"0000",
  7479 => x"0000",
  7480 => x"0000",
  7481 => x"0000",
  7482 => x"0000",
  7483 => x"0000",
  7484 => x"0000",
  7485 => x"0000",
  7486 => x"0000",
  7487 => x"0000",
  7488 => x"0000",
  7489 => x"0000",
  7490 => x"0000",
  7491 => x"0000",
  7492 => x"0000",
  7493 => x"0000",
  7494 => x"0000",
  7495 => x"0000",
  7496 => x"0000",
  7497 => x"0000",
  7498 => x"0000",
  7499 => x"0000",
  7500 => x"0000",
  7501 => x"0000",
  7502 => x"0000",
  7503 => x"0000",
  7504 => x"0000",
  7505 => x"0000",
  7506 => x"0000",
  7507 => x"0000",
  7508 => x"0000",
  7509 => x"0000",
  7510 => x"0000",
  7511 => x"0000",
  7512 => x"0000",
  7513 => x"0000",
  7514 => x"0000",
  7515 => x"0000",
  7516 => x"0000",
  7517 => x"0000",
  7518 => x"0000",
  7519 => x"0000",
  7520 => x"0000",
  7521 => x"0000",
  7522 => x"0000",
  7523 => x"0000",
  7524 => x"0000",
  7525 => x"0000",
  7526 => x"0000",
  7527 => x"0000",
  7528 => x"0000",
  7529 => x"0000",
  7530 => x"0000",
  7531 => x"0000",
  7532 => x"0000",
  7533 => x"0000",
  7534 => x"0000",
  7535 => x"0000",
  7536 => x"0000",
  7537 => x"0000",
  7538 => x"0000",
  7539 => x"0000",
  7540 => x"0000",
  7541 => x"0000",
  7542 => x"0000",
  7543 => x"0000",
  7544 => x"0000",
  7545 => x"0000",
  7546 => x"0000",
  7547 => x"0000",
  7548 => x"0000",
  7549 => x"0000",
  7550 => x"0000",
  7551 => x"0000",
  7552 => x"0000",
  7553 => x"0000",
  7554 => x"0000",
  7555 => x"0000",
  7556 => x"0000",
  7557 => x"0000",
  7558 => x"0000",
  7559 => x"0000",
  7560 => x"0000",
  7561 => x"0000",
  7562 => x"0000",
  7563 => x"0000",
  7564 => x"0000",
  7565 => x"0000",
  7566 => x"0000",
  7567 => x"0000",
  7568 => x"0000",
  7569 => x"0000",
  7570 => x"0000",
  7571 => x"0000",
  7572 => x"0000",
  7573 => x"0000",
  7574 => x"0000",
  7575 => x"0000",
  7576 => x"0000",
  7577 => x"0000",
  7578 => x"0000",
  7579 => x"0000",
  7580 => x"0000",
  7581 => x"0000",
  7582 => x"0000",
  7583 => x"0000",
  7584 => x"0000",
  7585 => x"0000",
  7586 => x"0000",
  7587 => x"0000",
  7588 => x"0000",
  7589 => x"0000",
  7590 => x"0000",
  7591 => x"0000",
  7592 => x"0000",
  7593 => x"0000",
  7594 => x"0000",
  7595 => x"0000",
  7596 => x"0000",
  7597 => x"0000",
  7598 => x"0000",
  7599 => x"0000",
  7600 => x"0000",
  7601 => x"0000",
  7602 => x"0000",
  7603 => x"0000",
  7604 => x"0000",
  7605 => x"0000",
  7606 => x"0000",
  7607 => x"0000",
  7608 => x"0000",
  7609 => x"0000",
  7610 => x"0000",
  7611 => x"0000",
  7612 => x"0000",
  7613 => x"0000",
  7614 => x"0000",
  7615 => x"0000",
  7616 => x"0000",
  7617 => x"0000",
  7618 => x"0000",
  7619 => x"0000",
  7620 => x"0000",
  7621 => x"0000",
  7622 => x"0000",
  7623 => x"0000",
  7624 => x"0000",
  7625 => x"0000",
  7626 => x"0000",
  7627 => x"0000",
  7628 => x"0000",
  7629 => x"0000",
  7630 => x"0000",
  7631 => x"0000",
  7632 => x"0000",
  7633 => x"0000",
  7634 => x"0000",
  7635 => x"0000",
  7636 => x"0000",
  7637 => x"0000",
  7638 => x"0000",
  7639 => x"0000",
  7640 => x"0000",
  7641 => x"0000",
  7642 => x"0000",
  7643 => x"0000",
  7644 => x"0000",
  7645 => x"0000",
  7646 => x"0000",
  7647 => x"0000",
  7648 => x"0000",
  7649 => x"0000",
  7650 => x"0000",
  7651 => x"0000",
  7652 => x"0000",
  7653 => x"0000",
  7654 => x"0000",
  7655 => x"0000",
  7656 => x"0000",
  7657 => x"0000",
  7658 => x"0000",
  7659 => x"0000",
  7660 => x"0000",
  7661 => x"0000",
  7662 => x"0000",
  7663 => x"0000",
  7664 => x"0000",
  7665 => x"0000",
  7666 => x"0000",
  7667 => x"0000",
  7668 => x"0000",
  7669 => x"0000",
  7670 => x"0000",
  7671 => x"0000",
  7672 => x"0000",
  7673 => x"0000",
  7674 => x"0000",
  7675 => x"0000",
  7676 => x"0000",
  7677 => x"0000",
  7678 => x"0000",
  7679 => x"0000",
  7680 => x"0000",
  7681 => x"0000",
  7682 => x"0000",
  7683 => x"0000",
  7684 => x"0000",
  7685 => x"0000",
  7686 => x"0000",
  7687 => x"0000",
  7688 => x"0000",
  7689 => x"0000",
  7690 => x"0000",
  7691 => x"0000",
  7692 => x"0000",
  7693 => x"0000",
  7694 => x"0000",
  7695 => x"0000",
  7696 => x"0000",
  7697 => x"0000",
  7698 => x"0000",
  7699 => x"0000",
  7700 => x"0000",
  7701 => x"0000",
  7702 => x"0000",
  7703 => x"0000",
  7704 => x"0000",
  7705 => x"0000",
  7706 => x"0000",
  7707 => x"0000",
  7708 => x"0000",
  7709 => x"0000",
  7710 => x"0000",
  7711 => x"0000",
  7712 => x"0000",
  7713 => x"0000",
  7714 => x"0000",
  7715 => x"0000",
  7716 => x"0000",
  7717 => x"0000",
  7718 => x"0000",
  7719 => x"0000",
  7720 => x"0000",
  7721 => x"0000",
  7722 => x"0000",
  7723 => x"0000",
  7724 => x"0000",
  7725 => x"0000",
  7726 => x"0000",
  7727 => x"0000",
  7728 => x"0000",
  7729 => x"0000",
  7730 => x"0000",
  7731 => x"0000",
  7732 => x"0000",
  7733 => x"0000",
  7734 => x"0000",
  7735 => x"0000",
  7736 => x"0000",
  7737 => x"0000",
  7738 => x"0000",
  7739 => x"0000",
  7740 => x"0000",
  7741 => x"0000",
  7742 => x"0000",
  7743 => x"0000",
  7744 => x"0000",
  7745 => x"0000",
  7746 => x"0000",
  7747 => x"0000",
  7748 => x"0000",
  7749 => x"0000",
  7750 => x"0000",
  7751 => x"0000",
  7752 => x"0000",
  7753 => x"0000",
  7754 => x"0000",
  7755 => x"0000",
  7756 => x"0000",
  7757 => x"0000",
  7758 => x"0000",
  7759 => x"0000",
  7760 => x"0000",
  7761 => x"0000",
  7762 => x"0000",
  7763 => x"0000",
  7764 => x"0000",
  7765 => x"0000",
  7766 => x"0000",
  7767 => x"0000",
  7768 => x"0000",
  7769 => x"0000",
  7770 => x"0000",
  7771 => x"0000",
  7772 => x"0000",
  7773 => x"0000",
  7774 => x"0000",
  7775 => x"0000",
  7776 => x"0000",
  7777 => x"0000",
  7778 => x"0000",
  7779 => x"0000",
  7780 => x"0000",
  7781 => x"0000",
  7782 => x"0000",
  7783 => x"0000",
  7784 => x"0000",
  7785 => x"0000",
  7786 => x"0000",
  7787 => x"0000",
  7788 => x"0000",
  7789 => x"0000",
  7790 => x"0000",
  7791 => x"0000",
  7792 => x"0000",
  7793 => x"0000",
  7794 => x"0000",
  7795 => x"0000",
  7796 => x"0000",
  7797 => x"0000",
  7798 => x"0000",
  7799 => x"0000",
  7800 => x"0000",
  7801 => x"0000",
  7802 => x"0000",
  7803 => x"0000",
  7804 => x"0000",
  7805 => x"0000",
  7806 => x"0000",
  7807 => x"0000",
  7808 => x"0000",
  7809 => x"0000",
  7810 => x"0000",
  7811 => x"0000",
  7812 => x"0000",
  7813 => x"0000",
  7814 => x"0000",
  7815 => x"0000",
  7816 => x"0000",
  7817 => x"0000",
  7818 => x"0000",
  7819 => x"0000",
  7820 => x"0000",
  7821 => x"0000",
  7822 => x"0000",
  7823 => x"0000",
  7824 => x"0000",
  7825 => x"0000",
  7826 => x"0000",
  7827 => x"0000",
  7828 => x"0000",
  7829 => x"0000",
  7830 => x"0000",
  7831 => x"0000",
  7832 => x"0000",
  7833 => x"0000",
  7834 => x"0000",
  7835 => x"0000",
  7836 => x"0000",
  7837 => x"0000",
  7838 => x"0000",
  7839 => x"0000",
  7840 => x"0000",
  7841 => x"0000",
  7842 => x"0000",
  7843 => x"0000",
  7844 => x"0000",
  7845 => x"0000",
  7846 => x"0000",
  7847 => x"0000",
  7848 => x"0000",
  7849 => x"0000",
  7850 => x"0000",
  7851 => x"0000",
  7852 => x"0000",
  7853 => x"0000",
  7854 => x"0000",
  7855 => x"0000",
  7856 => x"0000",
  7857 => x"0000",
  7858 => x"0000",
  7859 => x"0000",
  7860 => x"0000",
  7861 => x"0000",
  7862 => x"0000",
  7863 => x"0000",
  7864 => x"0000",
  7865 => x"0000",
  7866 => x"0000",
  7867 => x"0000",
  7868 => x"0000",
  7869 => x"0000",
  7870 => x"0000",
  7871 => x"0000",
  7872 => x"0000",
  7873 => x"0000",
  7874 => x"0000",
  7875 => x"0000",
  7876 => x"0000",
  7877 => x"0000",
  7878 => x"0000",
  7879 => x"0000",
  7880 => x"0000",
  7881 => x"0000",
  7882 => x"0000",
  7883 => x"0000",
  7884 => x"0000",
  7885 => x"0000",
  7886 => x"0000",
  7887 => x"0000",
  7888 => x"0000",
  7889 => x"0000",
  7890 => x"0000",
  7891 => x"0000",
  7892 => x"0000",
  7893 => x"0000",
  7894 => x"0000",
  7895 => x"0000",
  7896 => x"0000",
  7897 => x"0000",
  7898 => x"0000",
  7899 => x"0000",
  7900 => x"0000",
  7901 => x"0000",
  7902 => x"0000",
  7903 => x"0000",
  7904 => x"0000",
  7905 => x"0000",
  7906 => x"0000",
  7907 => x"0000",
  7908 => x"0000",
  7909 => x"0000",
  7910 => x"0000",
  7911 => x"0000",
  7912 => x"0000",
  7913 => x"0000",
  7914 => x"0000",
  7915 => x"0000",
  7916 => x"0000",
  7917 => x"0000",
  7918 => x"0000",
  7919 => x"0000",
  7920 => x"0000",
  7921 => x"0000",
  7922 => x"0000",
  7923 => x"0000",
  7924 => x"0000",
  7925 => x"0000",
  7926 => x"0000",
  7927 => x"0000",
  7928 => x"0000",
  7929 => x"0000",
  7930 => x"0000",
  7931 => x"0000",
  7932 => x"0000",
  7933 => x"0000",
  7934 => x"0000",
  7935 => x"0000",
  7936 => x"0000",
  7937 => x"0000",
  7938 => x"0000",
  7939 => x"0000",
  7940 => x"0000",
  7941 => x"0000",
  7942 => x"0000",
  7943 => x"0000",
  7944 => x"0000",
  7945 => x"0000",
  7946 => x"0000",
  7947 => x"0000",
  7948 => x"0000",
  7949 => x"0000",
  7950 => x"0000",
  7951 => x"0000",
  7952 => x"0000",
  7953 => x"0000",
  7954 => x"0000",
  7955 => x"0000",
  7956 => x"0000",
  7957 => x"0000",
  7958 => x"0000",
  7959 => x"0000",
  7960 => x"0000",
  7961 => x"0000",
  7962 => x"0000",
  7963 => x"0000",
  7964 => x"0000",
  7965 => x"0000",
  7966 => x"0000",
  7967 => x"0000",
  7968 => x"0000",
  7969 => x"0000",
  7970 => x"0000",
  7971 => x"0000",
  7972 => x"0000",
  7973 => x"0000",
  7974 => x"0000",
  7975 => x"0000",
  7976 => x"0000",
  7977 => x"0000",
  7978 => x"0000",
  7979 => x"0000",
  7980 => x"0000",
  7981 => x"0000",
  7982 => x"0000",
  7983 => x"0000",
  7984 => x"0000",
  7985 => x"0000",
  7986 => x"0000",
  7987 => x"0000",
  7988 => x"0000",
  7989 => x"0000",
  7990 => x"0000",
  7991 => x"0000",
  7992 => x"0000",
  7993 => x"0000",
  7994 => x"0000",
  7995 => x"0000",
  7996 => x"0000",
  7997 => x"0000",
  7998 => x"0000",
  7999 => x"0000",
  8000 => x"0000",
  8001 => x"0000",
  8002 => x"0000",
  8003 => x"0000",
  8004 => x"0000",
  8005 => x"0000",
  8006 => x"0000",
  8007 => x"0000",
  8008 => x"0000",
  8009 => x"0000",
  8010 => x"0000",
  8011 => x"0000",
  8012 => x"0000",
  8013 => x"0000",
  8014 => x"0000",
  8015 => x"0000",
  8016 => x"0000",
  8017 => x"0000",
  8018 => x"0000",
  8019 => x"0000",
  8020 => x"0000",
  8021 => x"0000",
  8022 => x"0000",
  8023 => x"0000",
  8024 => x"0000",
  8025 => x"0000",
  8026 => x"0000",
  8027 => x"0000",
  8028 => x"0000",
  8029 => x"0000",
  8030 => x"0000",
  8031 => x"0000",
  8032 => x"0000",
  8033 => x"0000",
  8034 => x"0000",
  8035 => x"0000",
  8036 => x"0000",
  8037 => x"0000",
  8038 => x"0000",
  8039 => x"0000",
  8040 => x"0000",
  8041 => x"0000",
  8042 => x"0000",
  8043 => x"0000",
  8044 => x"0000",
  8045 => x"0000",
  8046 => x"0000",
  8047 => x"0000",
  8048 => x"0000",
  8049 => x"0000",
  8050 => x"0000",
  8051 => x"0000",
  8052 => x"0000",
  8053 => x"0000",
  8054 => x"0000",
  8055 => x"0000",
  8056 => x"0000",
  8057 => x"0000",
  8058 => x"0000",
  8059 => x"0000",
  8060 => x"0000",
  8061 => x"0000",
  8062 => x"0000",
  8063 => x"0000",
  8064 => x"0000",
  8065 => x"0000",
  8066 => x"0000",
  8067 => x"0000",
  8068 => x"0000",
  8069 => x"0000",
  8070 => x"0000",
  8071 => x"0000",
  8072 => x"0000",
  8073 => x"0000",
  8074 => x"0000",
  8075 => x"0000",
  8076 => x"0000",
  8077 => x"0000",
  8078 => x"0000",
  8079 => x"0000",
  8080 => x"0000",
  8081 => x"0000",
  8082 => x"0000",
  8083 => x"0000",
  8084 => x"0000",
  8085 => x"0000",
  8086 => x"0000",
  8087 => x"0000",
  8088 => x"0000",
  8089 => x"0000",
  8090 => x"0000",
  8091 => x"0000",
  8092 => x"0000",
  8093 => x"0000",
  8094 => x"0000",
  8095 => x"0000",
  8096 => x"0000",
  8097 => x"0000",
  8098 => x"0000",
  8099 => x"0000",
  8100 => x"0000",
  8101 => x"0000",
  8102 => x"0000",
  8103 => x"0000",
  8104 => x"0000",
  8105 => x"0000",
  8106 => x"0000",
  8107 => x"0000",
  8108 => x"0000",
  8109 => x"0000",
  8110 => x"0000",
  8111 => x"0000",
  8112 => x"0000",
  8113 => x"0000",
  8114 => x"0000",
  8115 => x"0000",
  8116 => x"0000",
  8117 => x"0000",
  8118 => x"0000",
  8119 => x"0000",
  8120 => x"0000",
  8121 => x"0000",
  8122 => x"0000",
  8123 => x"0000",
  8124 => x"0000",
  8125 => x"0000",
  8126 => x"0000",
  8127 => x"0000",
  8128 => x"0000",
  8129 => x"0000",
  8130 => x"0000",
  8131 => x"0000",
  8132 => x"0000",
  8133 => x"0000",
  8134 => x"0000",
  8135 => x"0000",
  8136 => x"0000",
  8137 => x"0000",
  8138 => x"0000",
  8139 => x"0000",
  8140 => x"0000",
  8141 => x"0000",
  8142 => x"0000",
  8143 => x"0000",
  8144 => x"0000",
  8145 => x"0000",
  8146 => x"0000",
  8147 => x"0000",
  8148 => x"0000",
  8149 => x"0000",
  8150 => x"0000",
  8151 => x"0000",
  8152 => x"0000",
  8153 => x"0000",
  8154 => x"0000",
  8155 => x"0000",
  8156 => x"0000",
  8157 => x"0000",
  8158 => x"0000",
  8159 => x"0000",
  8160 => x"0000",
  8161 => x"0000",
  8162 => x"0000",
  8163 => x"0000",
  8164 => x"0000",
  8165 => x"0000",
  8166 => x"0000",
  8167 => x"0000",
  8168 => x"0000",
  8169 => x"0000",
  8170 => x"0000",
  8171 => x"0000",
  8172 => x"0000",
  8173 => x"0000",
  8174 => x"0000",
  8175 => x"0000",
  8176 => x"0000",
  8177 => x"0000",
  8178 => x"0000",
  8179 => x"0000",
  8180 => x"0000",
  8181 => x"0000",
  8182 => x"0000",
  8183 => x"0000",
  8184 => x"0000",
  8185 => x"0000",
  8186 => x"0000",
  8187 => x"0000",
  8188 => x"0000",
  8189 => x"0000",
  8190 => x"0000",
  8191 => x"0000",
  others => x"0000"
 );
begin
   process(CLK)
	begin 
		if (CLK'event AND CLK='1') then
			DOUT2 <= memoire(to_integer(unsigned(AD2)));
		end if;
	end process;

	process(CLK)
	begin 
		if (CLK'event AND CLK='1') then
			if ((CE1='1') AND (OE1='1')) then 
				DOUT1<=memoire(to_integer(unsigned(AD1)));
			else 
				DOUT1<=(others =>'0');
			end if;		
		end if;
	end process;
	
	process (CLK)
	begin
	  IF (CLK'event AND CLK='1') then
			if ((CE1='1') AND (WE1='1')) then 
				memoire(to_integer(unsigned(AD1)))<=DIN1;
			end if;
		  end if;
	end process;
	
end Behavioral;
