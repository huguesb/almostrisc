----------------------------------------------------------------------------------
--
-- File retrieved, on 07/02/2010, from :
-- http://sebastien-viardot.imag.fr/Enseignements/Archi1A2s/sources/ROMPROG.vhd
--
-- Slightly altered to get rid of vendor-specific packages and adjust formatting
-- Now auto-filled by asrom script
--
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROMPROG is
  Port ( AD : in  STD_LOGIC_VECTOR (12 downto 0);
         D : out  STD_LOGIC_VECTOR (15 downto 0);
         CLK : in STD_LOGIC);
end ROMPROG;

architecture Behavioral of ROMPROG is
  constant low_address: natural := 0;
  constant high_address: natural := 8192;
  subtype octet is std_logic_vector( 15 downto 0 );
  type zone_memoire is
    array (natural range low_address to high_address-1) of octet;
  constant m: zone_memoire:= (
    0=>x"FFF7",	-- 1111111111110111  liw	r7, IRQ_mask
    1=>x"2000",	-- 0010000000000000  
    2=>x"F8C0",	-- 1111100011000000  bai	-, os_init
    3=>x"0100",	-- 0000000100000000  
   16=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_ack
   17=>x"2002",	-- 0010000000000010  
   18=>x"D001",	-- 1101000000000001  lw	r1, r0
   19=>x"F54A",	-- 1111010101001010  bspl	r2, r1, 5
   20=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_error
   21=>x"0050",	-- 0000000001010000  
   22=>x"F4CA",	-- 1111010011001010  bspl	r2, r1, 3
   23=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_kbd
   24=>x"0060",	-- 0000000001100000  
   25=>x"F40A",	-- 1111010000001010  bspl	r2, r1, 0
   26=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_tmr
   27=>x"0040",	-- 0000000001000000  
   28=>x"D201",	-- 1101001000000001  sw	r1, r0
   29=>x"FFFE",	-- 1111111111111110  reti
   64=>x"263F",	-- 0010011000111111  not r7, r7
   65=>x"D7C0",	-- 1101011111000000  out	r7
   66=>x"E383",	-- 1110001110000011  ba	-, r6
   80=>x"25FF",	-- 0010010111111111  xor	r7, r7, r7
   81=>x"D7C0",	-- 1101011111000000  out	r7
   82=>x"E383",	-- 1110001110000011  ba	-, r6
   96=>x"FFF2",	-- 1111111111110010  liw	r2, PS2_rx
   97=>x"2004",	-- 0010000000000100  
   98=>x"D012",	-- 1101000000010010  lw	r2, r2
   99=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map + 8
  100=>x"1808",	-- 0001100000001000  
  101=>x"D01B",	-- 1101000000011011  lw	r3, r3
  102=>x"1EBF",	-- 0001111010111111  mixll	r7, r7, r2
  103=>x"C784",	-- 1100011110000100  li	r4, 0xF0
  104=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  105=>x"9760",	-- 1001011101100000  brieq	r4, int_kbd.release
  106=>x"C704",	-- 1100011100000100  li	r4, 0xE0
  107=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  108=>x"9520",	-- 1001010100100000  brieq	r4, int_kbd.extended
  109=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  110=>x"8B24",	-- 1000101100100100  brine	r4, int_kbd_ext
  111=>x"C3B4",	-- 1100001110110100  li	r4, 0x76
  112=>x"C044",	-- 1100000001000100  li	r4, 0x08
  113=>x"C31C",	-- 1100001100011100  li	r4, 0x63
  114=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  115=>x"80E4",	-- 1000000011100100  brine	r4, int_kbd_notup
  116=>x"C00D",	-- 1100000000001101  li	r5, 1
  117=>x"8E83",	-- 1000111010000011  bri	-, int_kbd_end
  118=>x"C30C",	-- 1100001100001100  li	r4, 0x61
  119=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  120=>x"80E4",	-- 1000000011100100  brine	r4, int_kbd_notleft
  121=>x"C015",	-- 1100000000010101  li	r5, 2
  122=>x"8D43",	-- 1000110101000011  bri	-, int_kbd_end
  123=>x"C304",	-- 1100001100000100  li	r4, 0x60
  124=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  125=>x"80E4",	-- 1000000011100100  brine	r4, int_kbd_notdown
  126=>x"C025",	-- 1100000000100101  li	r5, 4
  127=>x"8C03",	-- 1000110000000011  bri	-, int_kbd_end
  128=>x"C354",	-- 1100001101010100  li	r4, 0x6A
  129=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  130=>x"80E4",	-- 1000000011100100  brine	r4, int_kbd_notright
  131=>x"C045",	-- 1100000001000101  li	r5, 8
  132=>x"8AC3",	-- 1000101011000011  bri	-, int_kbd_end
  133=>x"C0EC",	-- 1100000011101100  li	r4, 0x1D
  134=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  135=>x"80E4",	-- 1000000011100100  brine	r4, int_kbd_notW
  136=>x"C00D",	-- 1100000000001101  li	r5, 1
  137=>x"8983",	-- 1000100110000011  bri	-, int_kbd_end
  138=>x"C0E4",	-- 1100000011100100  li	r4, 0x1C
  139=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  140=>x"80E4",	-- 1000000011100100  brine	r4, int_kbd_notA
  141=>x"C015",	-- 1100000000010101  li	r5, 2
  142=>x"8843",	-- 1000100001000011  bri	-, int_kbd_end
  143=>x"C0DC",	-- 1100000011011100  li	r4, 0x1B
  144=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  145=>x"80E4",	-- 1000000011100100  brine	r4, int_kbd_notS
  146=>x"C025",	-- 1100000000100101  li	r5, 4
  147=>x"8703",	-- 1000011100000011  bri	-, int_kbd_end
  148=>x"C11C",	-- 1100000100011100  li	r4, 0x23
  149=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  150=>x"80E4",	-- 1000000011100100  brine	r4, int_kbd_notD
  151=>x"C045",	-- 1100000001000101  li	r5, 8
  152=>x"85C3",	-- 1000010111000011  bri	-, int_kbd_end
  153=>x"8883",	-- 1000100010000011  bri	-, int_kbd_done
  154=>x"C3AC",	-- 1100001110101100  li	r4, 0x75
  155=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  156=>x"80E4",	-- 1000000011100100  brine	r4, int_kbd_ext_notup
  157=>x"C00D",	-- 1100000000001101  li	r5, 1
  158=>x"8443",	-- 1000010001000011  bri	-, int_kbd_end
  159=>x"C35C",	-- 1100001101011100  li	r4, 0x6B
  160=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  161=>x"80E4",	-- 1000000011100100  brine	r4, int_kbd_ext_notleft
  162=>x"C015",	-- 1100000000010101  li	r5, 2
  163=>x"8303",	-- 1000001100000011  bri	-, int_kbd_end
  164=>x"C394",	-- 1100001110010100  li	r4, 0x72
  165=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  166=>x"80E4",	-- 1000000011100100  brine	r4, int_kbd_ext_notdown
  167=>x"C025",	-- 1100000000100101  li	r5, 4
  168=>x"81C3",	-- 1000000111000011  bri	-, int_kbd_end
  169=>x"C3A4",	-- 1100001110100100  li	r4, 0x74
  170=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  171=>x"80E4",	-- 1000000011100100  brine	r4, int_kbd_ext_notright
  172=>x"C045",	-- 1100000001000101  li	r5, 8
  173=>x"8083",	-- 1000000010000011  bri	-, int_kbd_end
  174=>x"8343",	-- 1000001101000011  bri	-, int_kbd_done
  175=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  176=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  177=>x"1800",	-- 0001100000000000  
  178=>x"D01A",	-- 1101000000011010  lw	r2, r3
  179=>x"80E4",	-- 1000000011100100  brine	r4, int_kbd_maskout
  180=>x"2352",	-- 0010001101010010  or	r2, r2, r5
  181=>x"80C3",	-- 1000000011000011  bri	-, int_kbd_write
  182=>x"262D",	-- 0010011000101101  not	r5, r5
  183=>x"2152",	-- 0010000101010010  and	r2, r2, r5
  184=>x"D21A",	-- 1101001000011010  sw	r2, r3
  185=>x"C053",	-- 1100000001010011  li	r3, 10
  186=>x"D21A",	-- 1101001000011010  sw	r2, r3
  187=>x"C003",	-- 1100000000000011  li	r3, 0
  188=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  189=>x"1808",	-- 0001100000001000  
  190=>x"D223",	-- 1101001000100011  sw	r3, r4
  191=>x"E383",	-- 1110001110000011  ba	-, r6
  192=>x"C014",	-- 1100000000010100  li	r4, 2
  193=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  194=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  195=>x"1808",	-- 0001100000001000  
  196=>x"D223",	-- 1101001000100011  sw	r3, r4
  197=>x"E383",	-- 1110001110000011  ba	-, r6
  198=>x"C00C",	-- 1100000000001100  li	r4, 1
  199=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  200=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  201=>x"1808",	-- 0001100000001000  
  202=>x"D223",	-- 1101001000100011  sw	r3, r4
  203=>x"E383",	-- 1110001110000011  ba	-, r6
  256=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_mask
  257=>x"2000",	-- 0010000000000000  
  258=>x"C0C9",	-- 1100000011001001  li	r1, 0x19
  259=>x"D201",	-- 1101001000000001  sw	r1, r0
  260=>x"0400",	-- 0000010000000000  inc	r0, r0
  261=>x"CFF9",	-- 1100111111111001  li	r1, -1
  262=>x"D201",	-- 1101001000000001  sw	r1, r0
  263=>x"C03A",	-- 1100000000111010  li	r2, 7
  264=>x"0880",	-- 0000100010000000  add	r0, r0, r2
  265=>x"C0EA",	-- 1100000011101010  li	r2, 0x1D
  266=>x"D202",	-- 1101001000000010  sw	r2, r0
  267=>x"0400",	-- 0000010000000000  inc	r0, r0
  268=>x"C07A",	-- 1100000001111010  li	r2, 15
  269=>x"D202",	-- 1101001000000010  sw	r2, r0
  270=>x"FFF0",	-- 1111111111110000  liw	r0, key_press_map
  271=>x"1800",	-- 0001100000000000  
  272=>x"C001",	-- 1100000000000001  li	r1, 0
  273=>x"C042",	-- 1100000001000010  li	r2, 8
  274=>x"D201",	-- 1101001000000001  sw	r1, r0
  275=>x"0400",	-- 0000010000000000  inc	r0, r0
  276=>x"0612",	-- 0000011000010010  dec	r2, r2
  277=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  278=>x"C0F3",	-- 1100000011110011  li	r3, 30
  279=>x"CFFA",	-- 1100111111111010  li	r2, -1
  280=>x"D21A",	-- 1101001000011010  sw	r2, r3
  281=>x"8083",	-- 1000000010000011  bri	-, PaperGameStart
  282=>x"8003",	-- 1000000000000011  bri	-, PaperMenuLoop
  283=>x"FFF0",	-- 1111111111110000  liw	r0, paper_dir
  284=>x"1730",	-- 0001011100110000  
  285=>x"C001",	-- 1100000000000001  li	r1, 0
  286=>x"D201",	-- 1101001000000001  sw	r1, r0
  287=>x"0400",	-- 0000010000000000  inc	r0, r0
  288=>x"C4C1",	-- 1100010011000001  li	r1, 152
  289=>x"D201",	-- 1101001000000001  sw	r1, r0
  290=>x"0400",	-- 0000010000000000  inc	r0, r0
  291=>x"C001",	-- 1100000000000001  li	r1, 0
  292=>x"D201",	-- 1101001000000001  sw	r1, r0
  293=>x"0400",	-- 0000010000000000  inc	r0, r0
  294=>x"C401",	-- 1100010000000001  li	r1, 128
  295=>x"D201",	-- 1101001000000001  sw	r1, r0
  296=>x"0400",	-- 0000010000000000  inc	r0, r0
  297=>x"C001",	-- 1100000000000001  li	r1, 0
  298=>x"D201",	-- 1101001000000001  sw	r1, r0
  299=>x"0400",	-- 0000010000000000  inc	r0, r0
  300=>x"C0A1",	-- 1100000010100001  li	r1, 20
  301=>x"D201",	-- 1101001000000001  sw	r1, r0
  302=>x"0400",	-- 0000010000000000  inc	r0, r0
  303=>x"C029",	-- 1100000000101001  li	r1, 5
  304=>x"D201",	-- 1101001000000001  sw	r1, r0
  305=>x"0400",	-- 0000010000000000  inc	r0, r0
  306=>x"C000",	-- 1100000000000000  li	r0, 0
  307=>x"CFF9",	-- 1100111111111001  li	r1, -1
  308=>x"C0A2",	-- 1100000010100010  li	r2, 20
  309=>x"D201",	-- 1101001000000001  sw	r1, r0
  310=>x"0400",	-- 0000010000000000  inc	r0, r0
  311=>x"0612",	-- 0000011000010010  dec	r2, r2
  312=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  313=>x"C001",	-- 1100000000000001  li	r1, 0
  314=>x"FFF2",	-- 1111111111110010  liw	r2, 18*20
  315=>x"0168",	-- 0000000101101000  
  316=>x"D201",	-- 1101001000000001  sw	r1, r0
  317=>x"0400",	-- 0000010000000000  inc	r0, r0
  318=>x"0612",	-- 0000011000010010  dec	r2, r2
  319=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  320=>x"CFF9",	-- 1100111111111001  li	r1, -1
  321=>x"C0A2",	-- 1100000010100010  li	r2, 20
  322=>x"D201",	-- 1101001000000001  sw	r1, r0
  323=>x"0400",	-- 0000010000000000  inc	r0, r0
  324=>x"0612",	-- 0000011000010010  dec	r2, r2
  325=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  326=>x"C020",	-- 1100000000100000  li	r0, 4
  327=>x"C029",	-- 1100000000101001  li	r1, 5
  328=>x"FFF2",	-- 1111111111110010  liw	r2, paper_title
  329=>x"1738",	-- 0001011100111000  
  330=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  331=>x"01D1",	-- 0000000111010001  
  332=>x"C790",	-- 1100011110010000  li	r0, 242
  333=>x"C009",	-- 1100000000001001  li	r1, 1
  334=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud
  335=>x"1720",	-- 0001011100100000  
  336=>x"C043",	-- 1100000001000011  li	r3, 8
  337=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  338=>x"025C",	-- 0000001001011100  
  339=>x"C118",	-- 1100000100011000  li	r0, 35
  340=>x"C009",	-- 1100000000001001  li	r1, 1
  341=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  342=>x"173E",	-- 0001011100111110  
  343=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  344=>x"01D1",	-- 0000000111010001  
  345=>x"C790",	-- 1100011110010000  li	r0, 242
  346=>x"C051",	-- 1100000001010001  li	r1, 10
  347=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud + 4
  348=>x"1724",	-- 0001011100100100  
  349=>x"C043",	-- 1100000001000011  li	r3, 8
  350=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  351=>x"025C",	-- 0000001001011100  
  352=>x"C118",	-- 1100000100011000  li	r0, 35
  353=>x"C051",	-- 1100000001010001  li	r1, 10
  354=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  355=>x"173E",	-- 0001011100111110  
  356=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  357=>x"01D1",	-- 0000000111010001  
  358=>x"FFF0",	-- 1111111111110000  liw	r0, 20*20
  359=>x"0190",	-- 0000000110010000  
  360=>x"C001",	-- 1100000000000001  li	r1, 0
  361=>x"FFF2",	-- 1111111111110010  liw	r2, 220*20
  362=>x"1130",	-- 0001000100110000  
  363=>x"D201",	-- 1101001000000001  sw	r1, r0
  364=>x"0400",	-- 0000010000000000  inc	r0, r0
  365=>x"0612",	-- 0000011000010010  dec	r2, r2
  366=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  367=>x"FFF3",	-- 1111111111110011  liw	r3, paper_dir
  368=>x"1730",	-- 0001011100110000  
  369=>x"D01C",	-- 1101000000011100  lw	r4, r3
  370=>x"041B",	-- 0000010000011011  inc	r3, r3
  371=>x"D018",	-- 1101000000011000  lw	r0, r3
  372=>x"041B",	-- 0000010000011011  inc	r3, r3
  373=>x"FFF2",	-- 1111111111110010  liw	r2, paper_sprites
  374=>x"16D0",	-- 0001011011010000  
  375=>x"4624",	-- 0100011000100100  shl	r4, r4, 3
  376=>x"0912",	-- 0000100100010010  add	r2, r2, r4
  377=>x"C161",	-- 1100000101100001  li	r1, 44
  378=>x"C083",	-- 1100000010000011  li	r3, 16
  379=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_16
  380=>x"020C",	-- 0000001000001100  
  381=>x"FFF2",	-- 1111111111110010  liw	r2, paper_dir
  382=>x"1730",	-- 0001011100110000  
  383=>x"D010",	-- 1101000000010000  lw	r0, r2
  384=>x"0412",	-- 0000010000010010  inc	r2, r2
  385=>x"D011",	-- 1101000000010001  lw	r1, r2
  386=>x"0600",	-- 0000011000000000  dec	r0, r0
  387=>x"80C4",	-- 1000000011000100  brine	r0, $+3
  388=>x"0609",	-- 0000011000001001  dec	r1, r1
  389=>x"8103",	-- 1000000100000011  bri	-, $+4
  390=>x"0600",	-- 0000011000000000  dec	r0, r0
  391=>x"8084",	-- 1000000010000100  brine	r0, $+2
  392=>x"0409",	-- 0000010000001001  inc	r1, r1
  393=>x"D211",	-- 1101001000010001  sw	r1, r2
  394=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  395=>x"1800",	-- 0001100000000000  
  396=>x"D01B",	-- 1101000000011011  lw	r3, r3
  397=>x"BC18",	-- 1011110000011000  brieq	r3, PaperGameLoop
  398=>x"F7DC",	-- 1111011111011100  bspl	r4, r3, 15
  399=>x"84A0",	-- 1000010010100000  brieq	r4, PaperGameQuit
  400=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  401=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveUp
  402=>x"F49C",	-- 1111010010011100  bspl	r4, r3, 2
  403=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveDOWN
  404=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  405=>x"8160",	-- 1000000101100000  brieq	r4, PaperNoMoveLEFT
  406=>x"FFF2",	-- 1111111111110010  liw	r2, paper_dir
  407=>x"1730",	-- 0001011100110000  
  408=>x"C010",	-- 1100000000010000  li	r0, 2
  409=>x"D210",	-- 1101001000010000  sw	r0, r2
  410=>x"F4DC",	-- 1111010011011100  bspl	r4, r3, 3
  411=>x"8160",	-- 1000000101100000  brieq	r4, PaperNoMoveRIGHT
  412=>x"FFF2",	-- 1111111111110010  liw	r2, paper_dir
  413=>x"1730",	-- 0001011100110000  
  414=>x"C008",	-- 1100000000001000  li	r0, 1
  415=>x"D210",	-- 1101001000010000  sw	r0, r2
  416=>x"B183",	-- 1011000110000011  bri	-, PaperGameRedrawContent
  417=>x"FFFF",	-- 1111111111111111  reset
  418=>x"C750",	-- 1100011101010000  li	r0, 234
  419=>x"C1C2",	-- 1100000111000010  li	r2, 56
  420=>x"FAC6",	-- 1111101011000110  bail	-, r6, div_16_16
  421=>x"01BA",	-- 0000000110111010  
  422=>x"C448",	-- 1100010001001000  li	r0, 137
  423=>x"C472",	-- 1100010001110010  li	r2, 142
  424=>x"FAC6",	-- 1111101011000110  bail	-, r6, mult_16_16
  425=>x"01AE",	-- 0000000110101110  
  426=>x"C03A",	-- 1100000000111010  li r2, 7
  427=>x"FAC6",	-- 1111101011000110  bail	-, r6, fact_16
  428=>x"01C5",	-- 0000000111000101  
  429=>x"FFFF",	-- 1111111111111111  reset
  430=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  431=>x"2524",	-- 0010010100100100  xor	r4, r4, r4
  432=>x"C085",	-- 1100000010000101  li	r5, 16
  433=>x"0849",	-- 0000100001001001  add	r1, r1, r1
  434=>x"0C00",	-- 0000110000000000  adc	r0, r0, r0
  435=>x"0EDB",	-- 0000111011011011  sbc	r3, r3, r3
  436=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  437=>x"08C9",	-- 0000100011001001  add	r1, r1, r3
  438=>x"0D00",	-- 0000110100000000  adc	r0, r0, r4
  439=>x"062D",	-- 0000011000101101  dec	r5, r5
  440=>x"BE6C",	-- 1011111001101100  brine	r5, mult_16_16.loop
  441=>x"E383",	-- 1110001110000011  ba	-, r6
  442=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  443=>x"C084",	-- 1100000010000100  li	r4, 16
  444=>x"0800",	-- 0000100000000000  add	r0, r0, r0
  445=>x"0C49",	-- 0000110001001001  adc	r1, r1, r1
  446=>x"0A8B",	-- 0000101010001011  sub	r3, r1, r2
  447=>x"80DD",	-- 1000000011011101  brilt	r3, div_16_16.skip
  448=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  449=>x"0400",	-- 0000010000000000  inc	r0, r0
  450=>x"0624",	-- 0000011000100100  dec	r4, r4
  451=>x"BE64",	-- 1011111001100100  brine	r4, div_16_16.loop
  452=>x"E383",	-- 1110001110000011  ba	-, r6
  453=>x"2400",	-- 0010010000000000  xor	r0, r0, r0
  454=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  455=>x"8250",	-- 1000001001010000  brieq	r2, fact_16.end
  456=>x"0409",	-- 0000010000001001  inc	r1, r1
  457=>x"1008",	-- 0001000000001000  mova	r0, r1
  458=>x"FAC6",	-- 1111101011000110  bail	-, r6, mult_16_16
  459=>x"01AE",	-- 0000000110101110  
  460=>x"8104",	-- 1000000100000100  brine	r0, fact_16.overflow
  461=>x"01AE",	-- 0000000110101110  
  462=>x"0612",	-- 0000011000010010  dec	r2, r2
  463=>x"BE94",	-- 1011111010010100  brine	r2, fact_16.loop
  464=>x"E383",	-- 1110001110000011  ba	-, r6
  465=>x"063F",	-- 0000011000111111  dec	r7, r7
  466=>x"D23E",	-- 1101001000111110  sw	r6, r7
  467=>x"D013",	-- 1101000000010011  lw	r3, r2
  468=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  469=>x"84D8",	-- 1000010011011000  brieq	r3, puts.end
  470=>x"063F",	-- 0000011000111111  dec	r7, r7
  471=>x"D23A",	-- 1101001000111010  sw	r2, r7
  472=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  473=>x"01EB",	-- 0000000111101011  
  474=>x"D03A",	-- 1101000000111010  lw	r2, r7
  475=>x"043F",	-- 0000010000111111  inc	r7, r7
  476=>x"D013",	-- 1101000000010011  lw	r3, r2
  477=>x"4E1B",	-- 0100111000011011  shl	r3, r3, 7
  478=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  479=>x"8258",	-- 1000001001011000  brieq	r3, puts.end
  480=>x"063F",	-- 0000011000111111  dec	r7, r7
  481=>x"D23A",	-- 1101001000111010  sw	r2, r7
  482=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  483=>x"01EB",	-- 0000000111101011  
  484=>x"D03A",	-- 1101000000111010  lw	r2, r7
  485=>x"043F",	-- 0000010000111111  inc	r7, r7
  486=>x"0412",	-- 0000010000010010  inc	r2, r2
  487=>x"BB03",	-- 1011101100000011  bri	-, puts.loop
  488=>x"D03E",	-- 1101000000111110  lw	r6, r7
  489=>x"043F",	-- 0000010000111111  inc	r7, r7
  490=>x"E383",	-- 1110001110000011  ba	-, r6
  491=>x"063F",	-- 0000011000111111  dec	r7, r7
  492=>x"D23E",	-- 1101001000111110  sw	r6, r7
  493=>x"063F",	-- 0000011000111111  dec	r7, r7
  494=>x"D238",	-- 1101001000111000  sw	r0, r7
  495=>x"063F",	-- 0000011000111111  dec	r7, r7
  496=>x"D239",	-- 1101001000111001  sw	r1, r7
  497=>x"FFF2",	-- 1111111111110010  liw	r2, font_map
  498=>x"12C0",	-- 0001001011000000  
  499=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  500=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  501=>x"C043",	-- 1100000001000011  li	r3, 8
  502=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  503=>x"0236",	-- 0000001000110110  
  504=>x"D039",	-- 1101000000111001  lw	r1, r7
  505=>x"043F",	-- 0000010000111111  inc	r7, r7
  506=>x"D038",	-- 1101000000111000  lw	r0, r7
  507=>x"043F",	-- 0000010000111111  inc	r7, r7
  508=>x"0400",	-- 0000010000000000  inc	r0, r0
  509=>x"D03E",	-- 1101000000111110  lw	r6, r7
  510=>x"043F",	-- 0000010000111111  inc	r7, r7
  511=>x"E383",	-- 1110001110000011  ba	-, r6
  512=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  513=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  514=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  515=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  516=>x"C0A0",	-- 1100000010100000  li	r0, 20
  517=>x"D011",	-- 1101000000010001  lw	r1, r2
  518=>x"D221",	-- 1101001000100001  sw	r1, r4
  519=>x"0412",	-- 0000010000010010  inc	r2, r2
  520=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  521=>x"061B",	-- 0000011000011011  dec	r3, r3
  522=>x"BEDC",	-- 1011111011011100  brine	r3, put_sprite_16_aligned.loop
  523=>x"E383",	-- 1110001110000011  ba	-, r6
  524=>x"C07D",	-- 1100000001111101  li	r5, 15
  525=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  526=>x"6600",	-- 0110011000000000  shr	r0, r0, 3
  527=>x"BC68",	-- 1011110001101000  brieq	r5, put_sprite_16_aligned
  528=>x"062D",	-- 0000011000101101  dec	r5, r5
  529=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  530=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  531=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  532=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  533=>x"063F",	-- 0000011000111111  dec	r7, r7
  534=>x"D23B",	-- 1101001000111011  sw	r3, r7
  535=>x"D011",	-- 1101000000010001  lw	r1, r2
  536=>x"CFF8",	-- 1100111111111000  li	r0, -1
  537=>x"3D40",	-- 0011110101000000  rsr	r0, r0, r5
  538=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  539=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  540=>x"D023",	-- 1101000000100011  lw	r3, r4
  541=>x"2600",	-- 0010011000000000  not	r0, r0
  542=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  543=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  544=>x"D221",	-- 1101001000100001  sw	r1, r4
  545=>x"0424",	-- 0000010000100100  inc	r4, r4
  546=>x"D011",	-- 1101000000010001  lw	r1, r2
  547=>x"262D",	-- 0010011000101101  not	r5, r5
  548=>x"CFF8",	-- 1100111111111000  li	r0, -1
  549=>x"3F40",	-- 0011111101000000  rsl	r0, r0, r5
  550=>x"3B49",	-- 0011101101001001  rrl	r1, r1, r5
  551=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  552=>x"262D",	-- 0010011000101101  not	r5, r5
  553=>x"D023",	-- 1101000000100011  lw	r3, r4
  554=>x"2600",	-- 0010011000000000  not	r0, r0
  555=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  556=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  557=>x"D221",	-- 1101001000100001  sw	r1, r4
  558=>x"0412",	-- 0000010000010010  inc	r2, r2
  559=>x"C098",	-- 1100000010011000  li	r0, 19
  560=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  561=>x"D03B",	-- 1101000000111011  lw	r3, r7
  562=>x"043F",	-- 0000010000111111  inc	r7, r7
  563=>x"061B",	-- 0000011000011011  dec	r3, r3
  564=>x"B85C",	-- 1011100001011100  brine	r3, put_sprite_16.loop
  565=>x"E383",	-- 1110001110000011  ba	-, r6
  566=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  567=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  568=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  569=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  570=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  571=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  572=>x"C0A5",	-- 1100000010100101  li	r5, 20
  573=>x"8404",	-- 1000010000000100  brine	r0, put_sprite_8_aligned.loop1
  574=>x"D010",	-- 1101000000010000  lw	r0, r2
  575=>x"D021",	-- 1101000000100001  lw	r1, r4
  576=>x"1A41",	-- 0001101001000001  mixhl	r1, r0, r1
  577=>x"D221",	-- 1101001000100001  sw	r1, r4
  578=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  579=>x"061B",	-- 0000011000011011  dec	r3, r3
  580=>x"E398",	-- 1110001110011000  baeq	r3, r6
  581=>x"D021",	-- 1101000000100001  lw	r1, r4
  582=>x"1E41",	-- 0001111001000001  mixll	r1, r0, r1
  583=>x"D221",	-- 1101001000100001  sw	r1, r4
  584=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  585=>x"0412",	-- 0000010000010010  inc	r2, r2
  586=>x"061B",	-- 0000011000011011  dec	r3, r3
  587=>x"E398",	-- 1110001110011000  baeq	r3, r6
  588=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop0
  589=>x"D010",	-- 1101000000010000  lw	r0, r2
  590=>x"D021",	-- 1101000000100001  lw	r1, r4
  591=>x"1809",	-- 0001100000001001  mixhh	r1, r1, r0
  592=>x"D221",	-- 1101001000100001  sw	r1, r4
  593=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  594=>x"061B",	-- 0000011000011011  dec	r3, r3
  595=>x"E398",	-- 1110001110011000  baeq	r3, r6
  596=>x"D021",	-- 1101000000100001  lw	r1, r4
  597=>x"1A09",	-- 0001101000001001  mixhl	r1, r1, r0
  598=>x"D221",	-- 1101001000100001  sw	r1, r4
  599=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  600=>x"0412",	-- 0000010000010010  inc	r2, r2
  601=>x"061B",	-- 0000011000011011  dec	r3, r3
  602=>x"E398",	-- 1110001110011000  baeq	r3, r6
  603=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop1
  604=>x"C03D",	-- 1100000000111101  li	r5, 7
  605=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  606=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  607=>x"B5E8",	-- 1011010111101000  brieq	r5, put_sprite_8_aligned
  608=>x"062D",	-- 0000011000101101  dec	r5, r5
  609=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  610=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  611=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  612=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  613=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  614=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  615=>x"8A04",	-- 1000101000000100  brine	r0, put_sprite_8.loop1
  616=>x"D010",	-- 1101000000010000  lw	r0, r2
  617=>x"063F",	-- 0000011000111111  dec	r7, r7
  618=>x"D23A",	-- 1101001000111010  sw	r2, r7
  619=>x"C802",	-- 1100100000000010  li	r2, 0x100
  620=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  621=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  622=>x"D021",	-- 1101000000100001  lw	r1, r4
  623=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  624=>x"2612",	-- 0010011000010010  not	r2, r2
  625=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  626=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  627=>x"D221",	-- 1101001000100001  sw	r1, r4
  628=>x"C0A1",	-- 1100000010100001  li	r1, 20
  629=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  630=>x"D03A",	-- 1101000000111010  lw	r2, r7
  631=>x"043F",	-- 0000010000111111  inc	r7, r7
  632=>x"061B",	-- 0000011000011011  dec	r3, r3
  633=>x"E398",	-- 1110001110011000  baeq	r3, r6
  634=>x"D010",	-- 1101000000010000  lw	r0, r2
  635=>x"063F",	-- 0000011000111111  dec	r7, r7
  636=>x"D23A",	-- 1101001000111010  sw	r2, r7
  637=>x"1E00",	-- 0001111000000000  mixll	r0, r0, r0
  638=>x"C802",	-- 1100100000000010  li	r2, 0x100
  639=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  640=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  641=>x"D021",	-- 1101000000100001  lw	r1, r4
  642=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  643=>x"2612",	-- 0010011000010010  not	r2, r2
  644=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  645=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  646=>x"D221",	-- 1101001000100001  sw	r1, r4
  647=>x"C0A1",	-- 1100000010100001  li	r1, 20
  648=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  649=>x"D03A",	-- 1101000000111010  lw	r2, r7
  650=>x"043F",	-- 0000010000111111  inc	r7, r7
  651=>x"0412",	-- 0000010000010010  inc	r2, r2
  652=>x"061B",	-- 0000011000011011  dec	r3, r3
  653=>x"E398",	-- 1110001110011000  baeq	r3, r6
  654=>x"B683",	-- 1011011010000011  bri	-, put_sprite_8.loop0
  655=>x"D010",	-- 1101000000010000  lw	r0, r2
  656=>x"063F",	-- 0000011000111111  dec	r7, r7
  657=>x"D23A",	-- 1101001000111010  sw	r2, r7
  658=>x"063F",	-- 0000011000111111  dec	r7, r7
  659=>x"D23B",	-- 1101001000111011  sw	r3, r7
  660=>x"C802",	-- 1100100000000010  li	r2, 0x100
  661=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  662=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  663=>x"2080",	-- 0010000010000000  and	r0, r0, r2
  664=>x"D021",	-- 1101000000100001  lw	r1, r4
  665=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
  666=>x"261B",	-- 0010011000011011  not	r3, r3
  667=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  668=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
  669=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  670=>x"D221",	-- 1101001000100001  sw	r1, r4
  671=>x"0424",	-- 0000010000100100  inc	r4, r4
  672=>x"D021",	-- 1101000000100001  lw	r1, r4
  673=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  674=>x"261B",	-- 0010011000011011  not	r3, r3
  675=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  676=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
  677=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  678=>x"D221",	-- 1101001000100001  sw	r1, r4
  679=>x"C099",	-- 1100000010011001  li	r1, 19
  680=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  681=>x"D03B",	-- 1101000000111011  lw	r3, r7
  682=>x"043F",	-- 0000010000111111  inc	r7, r7
  683=>x"D03A",	-- 1101000000111010  lw	r2, r7
  684=>x"043F",	-- 0000010000111111  inc	r7, r7
  685=>x"061B",	-- 0000011000011011  dec	r3, r3
  686=>x"E398",	-- 1110001110011000  baeq	r3, r6
  687=>x"D010",	-- 1101000000010000  lw	r0, r2
  688=>x"4E00",	-- 0100111000000000  shl	r0, r0, 7
  689=>x"063F",	-- 0000011000111111  dec	r7, r7
  690=>x"D23A",	-- 1101001000111010  sw	r2, r7
  691=>x"063F",	-- 0000011000111111  dec	r7, r7
  692=>x"D23B",	-- 1101001000111011  sw	r3, r7
  693=>x"C802",	-- 1100100000000010  li	r2, 0x100
  694=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  695=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  696=>x"2080",	-- 0010000010000000  and	r0, r0, r2
  697=>x"D021",	-- 1101000000100001  lw	r1, r4
  698=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
  699=>x"261B",	-- 0010011000011011  not	r3, r3
  700=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  701=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
  702=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  703=>x"D221",	-- 1101001000100001  sw	r1, r4
  704=>x"0424",	-- 0000010000100100  inc	r4, r4
  705=>x"D021",	-- 1101000000100001  lw	r1, r4
  706=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  707=>x"261B",	-- 0010011000011011  not	r3, r3
  708=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  709=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
  710=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  711=>x"D221",	-- 1101001000100001  sw	r1, r4
  712=>x"C099",	-- 1100000010011001  li	r1, 19
  713=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  714=>x"D03B",	-- 1101000000111011  lw	r3, r7
  715=>x"043F",	-- 0000010000111111  inc	r7, r7
  716=>x"D03A",	-- 1101000000111010  lw	r2, r7
  717=>x"043F",	-- 0000010000111111  inc	r7, r7
  718=>x"0412",	-- 0000010000010010  inc	r2, r2
  719=>x"061B",	-- 0000011000011011  dec	r3, r3
  720=>x"E398",	-- 1110001110011000  baeq	r3, r6
  721=>x"AF83",	-- 1010111110000011  bri	-, put_sprite_8.loop1
    others => x"0000"
    );
begin
  process(CLK)
  begin
    if (CLK'event AND CLK='1') then
      D <= m(to_integer(unsigned(AD)));
    end if;
  end process;
end Behavioral;
