----------------------------------------------------------------------------------
--
-- File retrieved, on 07/02/2010, from :
-- http://sebastien-viardot.imag.fr/Enseignements/Archi1A2s/sources/ROMPROG.vhd
--
-- Slightly altered to get rid of vendor-specific packages and adjust formatting
--
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROMPROG is
  Port ( AD : in  STD_LOGIC_VECTOR (12 downto 0);
         D : out  STD_LOGIC_VECTOR (15 downto 0);
         CLK : in STD_LOGIC);
end ROMPROG;

architecture Behavioral of ROMPROG is
  constant low_address: natural := 0;
  constant high_address: natural := 8192;
  subtype octet is std_logic_vector( 15 downto 0 );
  type zone_memoire is
    array (natural range low_address to high_address-1) of octet;
  constant m: zone_memoire:= (
    0=>x"FFF7",	-- 1111111111110111  liw	r7, IRQ_mask
    1=>x"2000",	-- 0010000000000000  
    2=>x"F8C0",	-- 1111100011000000  bai	-, os_init
    3=>x"0100",	-- 0000000100000000  
   16=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_ack
   17=>x"2002",	-- 0010000000000010  
   18=>x"CFF9",	-- 1100111111111001  li	r1, -1
   19=>x"D201",	-- 1101001000000001  sw	r1, r0
   20=>x"261B",	-- 0010011000011011  not r3, r3
   21=>x"D6C0",	-- 1101011011000000  out	r3
   22=>x"FFFE",	-- 1111111111111110  reti
  256=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_mask
  257=>x"2000",	-- 0010000000000000  
  258=>x"C009",	-- 1100000000001001  li	r1, 1
  259=>x"D201",	-- 1101001000000001  sw	r1, r0
  260=>x"0400",	-- 0000010000000000  inc	r0, r0
  261=>x"CFF9",	-- 1100111111111001  li	r1, -1
  262=>x"D201",	-- 1101001000000001  sw	r1, r0
  263=>x"C03A",	-- 1100000000111010  li	r2, 7
  264=>x"0880",	-- 0000100010000000  add	r0, r0, r2
  265=>x"C0EA",	-- 1100000011101010  li	r2, 0x1D
  266=>x"D202",	-- 1101001000000010  sw	r2, r0
  267=>x"0400",	-- 0000010000000000  inc	r0, r0
  268=>x"C02A",	-- 1100000000101010  li	r2, 5
  269=>x"D202",	-- 1101001000000010  sw	r2, r0
  270=>x"FFF0",	-- 1111111111110000  liw	r0, 0x8421
  271=>x"8421",	-- 1000010000100001  
  272=>x"FFF1",	-- 1111111111110001  liw	r1, 0x1234
  273=>x"1234",	-- 0001001000110100  
  274=>x"E408",	-- 1110010000001000  exw	r0, r1
  275=>x"E408",	-- 1110010000001000  exw	r0, r1
  276=>x"1842",	-- 0001100001000010  mixhh	r2, r0, r1
  277=>x"1A43",	-- 0001101001000011  mixhl	r3, r0, r1
  278=>x"1C44",	-- 0001110001000100  mixlh	r4, r0, r1
  279=>x"1E45",	-- 0001111001000101  mixll	r5, r0, r1
  280=>x"C01E",	-- 1100000000011110  li	r6, 3
  281=>x"3985",	-- 0011100110000101  rrr	r5, r0, r6
  282=>x"3B8D",	-- 0011101110001101  rrl	r5, r1, r6
  283=>x"3D95",	-- 0011110110010101  rsr	r5, r2, r6
  284=>x"3F9D",	-- 0011111110011101  rsl	r5, r3, r6
  285=>x"FC0E",	-- 1111110000001110  mul	r6, r1, r0
  286=>x"C028",	-- 1100000000101000  li	r0, 5
  287=>x"C151",	-- 1100000101010001  li	r1, 42
  288=>x"FFF2",	-- 1111111111110010  liw	r2, font_map + 0x23 * 4
  289=>x"134C",	-- 0001001101001100  
  290=>x"C043",	-- 1100000001000011  li	r3, 8
  291=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  292=>x"019E",	-- 0000000110011110  
  293=>x"C000",	-- 1100000000000000  li	r0, 0
  294=>x"C0A1",	-- 1100000010100001  li	r1, 20
  295=>x"FFF2",	-- 1111111111110010  liw	r2, hello_str
  296=>x"16C0",	-- 0001011011000000  
  297=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  298=>x"015B",	-- 0000000101011011  
  299=>x"FFFF",	-- 1111111111111111  reset
  300=>x"C750",	-- 1100011101010000  li	r0, 234
  301=>x"C1C2",	-- 1100000111000010  li	r2, 56
  302=>x"FAC6",	-- 1111101011000110  bail	-, r6, div_16_16
  303=>x"0144",	-- 0000000101000100  
  304=>x"C448",	-- 1100010001001000  li	r0, 137
  305=>x"C472",	-- 1100010001110010  li	r2, 142
  306=>x"FAC6",	-- 1111101011000110  bail	-, r6, mult_16_16
  307=>x"0138",	-- 0000000100111000  
  308=>x"C03A",	-- 1100000000111010  li r2, 7
  309=>x"FAC6",	-- 1111101011000110  bail	-, r6, fact_16
  310=>x"014F",	-- 0000000101001111  
  311=>x"FFFF",	-- 1111111111111111  reset
  312=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  313=>x"2524",	-- 0010010100100100  xor	r4, r4, r4
  314=>x"C085",	-- 1100000010000101  li	r5, 16
  315=>x"0849",	-- 0000100001001001  add	r1, r1, r1
  316=>x"0C00",	-- 0000110000000000  adc	r0, r0, r0
  317=>x"0EDB",	-- 0000111011011011  sbc	r3, r3, r3
  318=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  319=>x"08C9",	-- 0000100011001001  add	r1, r1, r3
  320=>x"0D00",	-- 0000110100000000  adc	r0, r0, r4
  321=>x"062D",	-- 0000011000101101  dec	r5, r5
  322=>x"BE6C",	-- 1011111001101100  brine	r5, mult_16_16.loop
  323=>x"E383",	-- 1110001110000011  ba	-, r6
  324=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  325=>x"C084",	-- 1100000010000100  li	r4, 16
  326=>x"0800",	-- 0000100000000000  add	r0, r0, r0
  327=>x"0C49",	-- 0000110001001001  adc	r1, r1, r1
  328=>x"0A8B",	-- 0000101010001011  sub	r3, r1, r2
  329=>x"80DD",	-- 1000000011011101  brilt	r3, div_16_16.skip
  330=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  331=>x"0400",	-- 0000010000000000  inc	r0, r0
  332=>x"0624",	-- 0000011000100100  dec	r4, r4
  333=>x"BE64",	-- 1011111001100100  brine	r4, div_16_16.loop
  334=>x"E383",	-- 1110001110000011  ba	-, r6
  335=>x"2400",	-- 0010010000000000  xor	r0, r0, r0
  336=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  337=>x"8250",	-- 1000001001010000  brieq	r2, fact_16.end
  338=>x"0409",	-- 0000010000001001  inc	r1, r1
  339=>x"1008",	-- 0001000000001000  mova	r0, r1
  340=>x"FAC6",	-- 1111101011000110  bail	-, r6, mult_16_16
  341=>x"0138",	-- 0000000100111000  
  342=>x"8104",	-- 1000000100000100  brine	r0, fact_16.overflow
  343=>x"0138",	-- 0000000100111000  
  344=>x"0612",	-- 0000011000010010  dec	r2, r2
  345=>x"BE94",	-- 1011111010010100  brine	r2, fact_16.loop
  346=>x"E383",	-- 1110001110000011  ba	-, r6
  347=>x"D013",	-- 1101000000010011  lw	r3, r2
  348=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  349=>x"E398",	-- 1110001110011000  baeq	r3, r6
  350=>x"063F",	-- 0000011000111111  dec	r7, r7
  351=>x"D23E",	-- 1101001000111110  sw	r6, r7
  352=>x"063F",	-- 0000011000111111  dec	r7, r7
  353=>x"D238",	-- 1101001000111000  sw	r0, r7
  354=>x"063F",	-- 0000011000111111  dec	r7, r7
  355=>x"D239",	-- 1101001000111001  sw	r1, r7
  356=>x"063F",	-- 0000011000111111  dec	r7, r7
  357=>x"D23A",	-- 1101001000111010  sw	r2, r7
  358=>x"FFF4",	-- 1111111111110100  liw	r4, font_map
  359=>x"12C0",	-- 0001001011000000  
  360=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  361=>x"091A",	-- 0000100100011010  add	r2, r3, r4
  362=>x"C043",	-- 1100000001000011  li	r3, 8
  363=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  364=>x"019E",	-- 0000000110011110  
  365=>x"D03A",	-- 1101000000111010  lw	r2, r7
  366=>x"043F",	-- 0000010000111111  inc	r7, r7
  367=>x"D039",	-- 1101000000111001  lw	r1, r7
  368=>x"043F",	-- 0000010000111111  inc	r7, r7
  369=>x"D038",	-- 1101000000111000  lw	r0, r7
  370=>x"043F",	-- 0000010000111111  inc	r7, r7
  371=>x"D03E",	-- 1101000000111110  lw	r6, r7
  372=>x"043F",	-- 0000010000111111  inc	r7, r7
  373=>x"0400",	-- 0000010000000000  inc	r0, r0
  374=>x"D013",	-- 1101000000010011  lw	r3, r2
  375=>x"4E1B",	-- 0100111000011011  shl	r3, r3, 7
  376=>x"6A1B",	-- 0110101000011011  shr	r3, r3, 5
  377=>x"E398",	-- 1110001110011000  baeq	r3, r6
  378=>x"063F",	-- 0000011000111111  dec	r7, r7
  379=>x"D23E",	-- 1101001000111110  sw	r6, r7
  380=>x"063F",	-- 0000011000111111  dec	r7, r7
  381=>x"D238",	-- 1101001000111000  sw	r0, r7
  382=>x"063F",	-- 0000011000111111  dec	r7, r7
  383=>x"D239",	-- 1101001000111001  sw	r1, r7
  384=>x"063F",	-- 0000011000111111  dec	r7, r7
  385=>x"D23A",	-- 1101001000111010  sw	r2, r7
  386=>x"FFF4",	-- 1111111111110100  liw	r4, font_map
  387=>x"12C0",	-- 0001001011000000  
  388=>x"091A",	-- 0000100100011010  add	r2, r3, r4
  389=>x"C043",	-- 1100000001000011  li	r3, 8
  390=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  391=>x"019E",	-- 0000000110011110  
  392=>x"D03A",	-- 1101000000111010  lw	r2, r7
  393=>x"043F",	-- 0000010000111111  inc	r7, r7
  394=>x"D039",	-- 1101000000111001  lw	r1, r7
  395=>x"043F",	-- 0000010000111111  inc	r7, r7
  396=>x"D038",	-- 1101000000111000  lw	r0, r7
  397=>x"043F",	-- 0000010000111111  inc	r7, r7
  398=>x"D03E",	-- 1101000000111110  lw	r6, r7
  399=>x"043F",	-- 0000010000111111  inc	r7, r7
  400=>x"0400",	-- 0000010000000000  inc	r0, r0
  401=>x"0412",	-- 0000010000010010  inc	r2, r2
  402=>x"B243",	-- 1011001001000011  bri	-, puts.loop
  403=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  404=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  405=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  406=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  407=>x"D011",	-- 1101000000010001  lw	r1, r2
  408=>x"D221",	-- 1101001000100001  sw	r1, r4
  409=>x"0412",	-- 0000010000010010  inc	r2, r2
  410=>x"0424",	-- 0000010000100100  inc	r4, r4
  411=>x"061B",	-- 0000011000011011  dec	r3, r3
  412=>x"BEDC",	-- 1011111011011100  brine	r3, put_sprite_16_aligned.loop
  413=>x"E383",	-- 1110001110000011  ba	-, r6
  414=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  415=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  416=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  417=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  418=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  419=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  420=>x"C0A5",	-- 1100000010100101  li	r5, 20
  421=>x"8404",	-- 1000010000000100  brine	r0, put_sprite_8_aligned.loop1
  422=>x"D010",	-- 1101000000010000  lw	r0, r2
  423=>x"D021",	-- 1101000000100001  lw	r1, r4
  424=>x"1A41",	-- 0001101001000001  mixhl	r1, r0, r1
  425=>x"D221",	-- 1101001000100001  sw	r1, r4
  426=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  427=>x"061B",	-- 0000011000011011  dec	r3, r3
  428=>x"E398",	-- 1110001110011000  baeq	r3, r6
  429=>x"D021",	-- 1101000000100001  lw	r1, r4
  430=>x"1E41",	-- 0001111001000001  mixll	r1, r0, r1
  431=>x"D221",	-- 1101001000100001  sw	r1, r4
  432=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  433=>x"0412",	-- 0000010000010010  inc	r2, r2
  434=>x"061B",	-- 0000011000011011  dec	r3, r3
  435=>x"E398",	-- 1110001110011000  baeq	r3, r6
  436=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop0
  437=>x"D010",	-- 1101000000010000  lw	r0, r2
  438=>x"D021",	-- 1101000000100001  lw	r1, r4
  439=>x"1809",	-- 0001100000001001  mixhh	r1, r1, r0
  440=>x"D221",	-- 1101001000100001  sw	r1, r4
  441=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  442=>x"061B",	-- 0000011000011011  dec	r3, r3
  443=>x"E398",	-- 1110001110011000  baeq	r3, r6
  444=>x"D021",	-- 1101000000100001  lw	r1, r4
  445=>x"1A09",	-- 0001101000001001  mixhl	r1, r1, r0
  446=>x"D221",	-- 1101001000100001  sw	r1, r4
  447=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  448=>x"0412",	-- 0000010000010010  inc	r2, r2
  449=>x"061B",	-- 0000011000011011  dec	r3, r3
  450=>x"E398",	-- 1110001110011000  baeq	r3, r6
  451=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop1
    others => x"0000"
    );
begin
  process(CLK)
  begin
    if (CLK'event AND CLK='1') then
      D <= m(to_integer(unsigned(AD)));
    end if;
  end process;
end Behavioral;
