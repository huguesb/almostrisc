----------------------------------------------------------------------------------
--
-- File retrieved, on 07/02/2010, from :
-- http://sebastien-viardot.imag.fr/Enseignements/Archi1A2s/sources/ROMPROG.vhd
--
-- Slightly altered to get rid of vendor-specific packages and adjust formatting
-- Now auto-filled by asrom script
--
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROMPROG is
  Port ( AD : in  STD_LOGIC_VECTOR (12 downto 0);
         D : out  STD_LOGIC_VECTOR (15 downto 0);
         CLK : in STD_LOGIC);
end ROMPROG;

architecture Behavioral of ROMPROG is
  constant low_address: natural := 0;
  constant high_address: natural := 8192;
  subtype octet is std_logic_vector( 15 downto 0 );
  type zone_memoire is
    array (natural range low_address to high_address-1) of octet;
  constant m: zone_memoire:= (
    0=>x"FFF7",	-- 1111111111110111  liw	r7, IRQ_mask
    1=>x"2000",	-- 0010000000000000  
    2=>x"F8C0",	-- 1111100011000000  bai	-, os_init
    3=>x"0100",	-- 0000000100000000  
   16=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_ack
   17=>x"2002",	-- 0010000000000010  
   18=>x"D001",	-- 1101000000000001  lw	r1, r0
   19=>x"F54A",	-- 1111010101001010  bspl	r2, r1, 5
   20=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_error
   21=>x"0050",	-- 0000000001010000  
   22=>x"F4CA",	-- 1111010011001010  bspl	r2, r1, 3
   23=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_kbd
   24=>x"0060",	-- 0000000001100000  
   25=>x"F40A",	-- 1111010000001010  bspl	r2, r1, 0
   26=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_tmr
   27=>x"0040",	-- 0000000001000000  
   28=>x"D201",	-- 1101001000000001  sw	r1, r0
   29=>x"FFFE",	-- 1111111111111110  reti
   64=>x"263F",	-- 0010011000111111  not r7, r7
   65=>x"D7C0",	-- 1101011111000000  out	r7
   66=>x"E383",	-- 1110001110000011  ba	-, r6
   80=>x"25FF",	-- 0010010111111111  xor	r7, r7, r7
   81=>x"D7C0",	-- 1101011111000000  out	r7
   82=>x"E383",	-- 1110001110000011  ba	-, r6
   96=>x"FFF2",	-- 1111111111110010  liw	r2, PS2_rx
   97=>x"2004",	-- 0010000000000100  
   98=>x"D012",	-- 1101000000010010  lw	r2, r2
   99=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map + 8
  100=>x"16C8",	-- 0001011011001000  
  101=>x"D01B",	-- 1101000000011011  lw	r3, r3
  102=>x"1EBF",	-- 0001111010111111  mixll	r7, r7, r2
  103=>x"C784",	-- 1100011110000100  li	r4, 0xF0
  104=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  105=>x"8C60",	-- 1000110001100000  brieq	r4, int_kbd.release
  106=>x"C704",	-- 1100011100000100  li	r4, 0xE0
  107=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  108=>x"8A20",	-- 1000101000100000  brieq	r4, int_kbd.extended
  109=>x"FFF5",	-- 1111111111110101  liw	r5, rand_seed
  110=>x"16C8",	-- 0001011011001000  
  111=>x"D02C",	-- 1101000000101100  lw	r4, r5
  112=>x"24A4",	-- 0010010010100100  xor	r4, r4, r2
  113=>x"D22C",	-- 1101001000101100  sw	r4, r5
  114=>x"FFF5",	-- 1111111111110101  liw	r5, paper_keys - 1
  115=>x"16CF",	-- 0001011011001111  
  116=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  117=>x"80E0",	-- 1000000011100000  brieq	r4, $+3
  118=>x"FFF5",	-- 1111111111110101  liw	r5, paper_keys + 11 - 1
  119=>x"16DA",	-- 0001011011011010  
  120=>x"042D",	-- 0000010000101101  inc	r5, r5
  121=>x"D02C",	-- 1101000000101100  lw	r4, r5
  122=>x"8560",	-- 1000010101100000  brieq	r4, scan_code_mismatch
  123=>x"6E24",	-- 0110111000100100  shr	r4, r4, 7
  124=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  125=>x"BEE4",	-- 1011111011100100  brine	r4, scan_code_loop
  126=>x"D02A",	-- 1101000000101010  lw	r2, r5
  127=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  128=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  129=>x"741B",	-- 0111010000011011  shr	r3, r3, 10
  130=>x"C00D",	-- 1100000000001101  li	r5, 1
  131=>x"0612",	-- 0000011000010010  dec	r2, r2
  132=>x"3AAA",	-- 0011101010101010  rrl	r2, r5, r2
  133=>x"FFF5",	-- 1111111111110101  liw	r5, key_press_map
  134=>x"16C0",	-- 0001011011000000  
  135=>x"08ED",	-- 0000100011101101  add	r5, r5, r3
  136=>x"D02B",	-- 1101000000101011  lw	r3, r5
  137=>x"80E4",	-- 1000000011100100  brine	r4, scan_code_release
  138=>x"229B",	-- 0010001010011011  or	r3, r3, r2
  139=>x"80C3",	-- 1000000011000011  bri	-, scan_code_notify
  140=>x"2612",	-- 0010011000010010  not	r2, r2
  141=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  142=>x"D22B",	-- 1101001000101011  sw	r3, r5
  143=>x"C003",	-- 1100000000000011  li	r3, 0
  144=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  145=>x"16C8",	-- 0001011011001000  
  146=>x"D223",	-- 1101001000100011  sw	r3, r4
  147=>x"E383",	-- 1110001110000011  ba	-, r6
  148=>x"C014",	-- 1100000000010100  li	r4, 2
  149=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  150=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  151=>x"16C8",	-- 0001011011001000  
  152=>x"D223",	-- 1101001000100011  sw	r3, r4
  153=>x"E383",	-- 1110001110000011  ba	-, r6
  154=>x"C00C",	-- 1100000000001100  li	r4, 1
  155=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  156=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  157=>x"16C8",	-- 0001011011001000  
  158=>x"D223",	-- 1101001000100011  sw	r3, r4
  159=>x"E383",	-- 1110001110000011  ba	-, r6
  256=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_mask
  257=>x"2000",	-- 0010000000000000  
  258=>x"C0C9",	-- 1100000011001001  li	r1, 0x19
  259=>x"D201",	-- 1101001000000001  sw	r1, r0
  260=>x"0400",	-- 0000010000000000  inc	r0, r0
  261=>x"CFF9",	-- 1100111111111001  li	r1, -1
  262=>x"D201",	-- 1101001000000001  sw	r1, r0
  263=>x"C03A",	-- 1100000000111010  li	r2, 7
  264=>x"0880",	-- 0000100010000000  add	r0, r0, r2
  265=>x"C0EA",	-- 1100000011101010  li	r2, 0x1D
  266=>x"D202",	-- 1101001000000010  sw	r2, r0
  267=>x"0400",	-- 0000010000000000  inc	r0, r0
  268=>x"C07A",	-- 1100000001111010  li	r2, 15
  269=>x"D202",	-- 1101001000000010  sw	r2, r0
  270=>x"0400",	-- 0000010000000000  inc	r0, r0
  271=>x"C0DA",	-- 1100000011011010  li	r2, 0x1B
  272=>x"D202",	-- 1101001000000010  sw	r2, r0
  273=>x"0400",	-- 0000010000000000  inc	r0, r0
  274=>x"FFF2",	-- 1111111111110010  liw	r2, 817
  275=>x"0331",	-- 0000001100110001  
  276=>x"D202",	-- 1101001000000010  sw	r2, r0
  277=>x"FFF0",	-- 1111111111110000  liw	r0, key_press_map
  278=>x"16C0",	-- 0001011011000000  
  279=>x"C001",	-- 1100000000000001  li	r1, 0
  280=>x"C042",	-- 1100000001000010  li	r2, 8
  281=>x"D201",	-- 1101001000000001  sw	r1, r0
  282=>x"0400",	-- 0000010000000000  inc	r0, r0
  283=>x"0612",	-- 0000011000010010  dec	r2, r2
  284=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  285=>x"8083",	-- 1000000010000011  bri	-, PaperGameStart
  286=>x"8003",	-- 1000000000000011  bri	-, PaperMenuLoop
  287=>x"FFF0",	-- 1111111111110000  liw	r0, paper_score
  288=>x"16C9",	-- 0001011011001001  
  289=>x"C001",	-- 1100000000000001  li	r1, 0
  290=>x"D201",	-- 1101001000000001  sw	r1, r0
  291=>x"FFF0",	-- 1111111111110000  liw	r0, paper_dir
  292=>x"179C",	-- 0001011110011100  
  293=>x"C001",	-- 1100000000000001  li	r1, 0
  294=>x"D201",	-- 1101001000000001  sw	r1, r0
  295=>x"0400",	-- 0000010000000000  inc	r0, r0
  296=>x"FFF1",	-- 1111111111110001  liw	r1, 152 * 8
  297=>x"04C0",	-- 0000010011000000  
  298=>x"D201",	-- 1101001000000001  sw	r1, r0
  299=>x"0400",	-- 0000010000000000  inc	r0, r0
  300=>x"C001",	-- 1100000000000001  li	r1, 0
  301=>x"D201",	-- 1101001000000001  sw	r1, r0
  302=>x"0400",	-- 0000010000000000  inc	r0, r0
  303=>x"FFF1",	-- 1111111111110001  liw	r1, 128 * 8
  304=>x"0400",	-- 0000010000000000  
  305=>x"D201",	-- 1101001000000001  sw	r1, r0
  306=>x"0400",	-- 0000010000000000  inc	r0, r0
  307=>x"C001",	-- 1100000000000001  li	r1, 0
  308=>x"D201",	-- 1101001000000001  sw	r1, r0
  309=>x"0400",	-- 0000010000000000  inc	r0, r0
  310=>x"C069",	-- 1100000001101001  li	r1, 13
  311=>x"D201",	-- 1101001000000001  sw	r1, r0
  312=>x"0400",	-- 0000010000000000  inc	r0, r0
  313=>x"C011",	-- 1100000000010001  li	r1, 2
  314=>x"D201",	-- 1101001000000001  sw	r1, r0
  315=>x"0400",	-- 0000010000000000  inc	r0, r0
  316=>x"FFF0",	-- 1111111111110000  liw	r0, paper_tilemap
  317=>x"17B0",	-- 0001011110110000  
  318=>x"C001",	-- 1100000000000001  li	r1, 0
  319=>x"C0C2",	-- 1100000011000010  li	r2, 6*4
  320=>x"D201",	-- 1101001000000001  sw	r1, r0
  321=>x"0400",	-- 0000010000000000  inc	r0, r0
  322=>x"0612",	-- 0000011000010010  dec	r2, r2
  323=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  324=>x"C000",	-- 1100000000000000  li	r0, 0
  325=>x"CFF9",	-- 1100111111111001  li	r1, -1
  326=>x"C0A2",	-- 1100000010100010  li	r2, 20
  327=>x"D201",	-- 1101001000000001  sw	r1, r0
  328=>x"0400",	-- 0000010000000000  inc	r0, r0
  329=>x"0612",	-- 0000011000010010  dec	r2, r2
  330=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  331=>x"C001",	-- 1100000000000001  li	r1, 0
  332=>x"FFF2",	-- 1111111111110010  liw	r2, 18*20
  333=>x"0168",	-- 0000000101101000  
  334=>x"D201",	-- 1101001000000001  sw	r1, r0
  335=>x"0400",	-- 0000010000000000  inc	r0, r0
  336=>x"0612",	-- 0000011000010010  dec	r2, r2
  337=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  338=>x"CFF9",	-- 1100111111111001  li	r1, -1
  339=>x"C0A2",	-- 1100000010100010  li	r2, 20
  340=>x"D201",	-- 1101001000000001  sw	r1, r0
  341=>x"0400",	-- 0000010000000000  inc	r0, r0
  342=>x"0612",	-- 0000011000010010  dec	r2, r2
  343=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  344=>x"C020",	-- 1100000000100000  li	r0, 4
  345=>x"C029",	-- 1100000000101001  li	r1, 5
  346=>x"FFF2",	-- 1111111111110010  liw	r2, paper_title
  347=>x"17A4",	-- 0001011110100100  
  348=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  349=>x"02BD",	-- 0000001010111101  
  350=>x"C090",	-- 1100000010010000  li	r0, 18
  351=>x"C029",	-- 1100000000101001  li	r1, 5
  352=>x"FFF2",	-- 1111111111110010  liw	r2, paper_score
  353=>x"16C9",	-- 0001011011001001  
  354=>x"D012",	-- 1101000000010010  lw	r2, r2
  355=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum
  356=>x"02EC",	-- 0000001011101100  
  357=>x"C778",	-- 1100011101111000  li	r0, 239
  358=>x"C009",	-- 1100000000001001  li	r1, 1
  359=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud
  360=>x"1780",	-- 0001011110000000  
  361=>x"C043",	-- 1100000001000011  li	r3, 8
  362=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  363=>x"03C5",	-- 0000001111000101  
  364=>x"C0F8",	-- 1100000011111000  li	r0, 31
  365=>x"C009",	-- 1100000000001001  li	r1, 1
  366=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  367=>x"17A0",	-- 0001011110100000  
  368=>x"D012",	-- 1101000000010010  lw	r2, r2
  369=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum
  370=>x"02EC",	-- 0000001011101100  
  371=>x"C120",	-- 1100000100100000  li	r0, 36
  372=>x"C009",	-- 1100000000001001  li	r1, 1
  373=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  374=>x"17AA",	-- 0001011110101010  
  375=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  376=>x"02BD",	-- 0000001010111101  
  377=>x"C778",	-- 1100011101111000  li	r0, 239
  378=>x"C051",	-- 1100000001010001  li	r1, 10
  379=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud + 8
  380=>x"1788",	-- 0001011110001000  
  381=>x"C043",	-- 1100000001000011  li	r3, 8
  382=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  383=>x"03C5",	-- 0000001111000101  
  384=>x"C0F8",	-- 1100000011111000  li	r0, 31
  385=>x"C051",	-- 1100000001010001  li	r1, 10
  386=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed + 1
  387=>x"17A1",	-- 0001011110100001  
  388=>x"D012",	-- 1101000000010010  lw	r2, r2
  389=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum
  390=>x"02EC",	-- 0000001011101100  
  391=>x"C120",	-- 1100000100100000  li	r0, 36
  392=>x"C051",	-- 1100000001010001  li	r1, 10
  393=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  394=>x"17AA",	-- 0001011110101010  
  395=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  396=>x"02BD",	-- 0000001010111101  
  397=>x"FFF0",	-- 1111111111110000  liw	r0, 20*20
  398=>x"0190",	-- 0000000110010000  
  399=>x"C001",	-- 1100000000000001  li	r1, 0
  400=>x"FFF2",	-- 1111111111110010  liw	r2, 220*20
  401=>x"1130",	-- 0001000100110000  
  402=>x"D201",	-- 1101001000000001  sw	r1, r0
  403=>x"0400",	-- 0000010000000000  inc	r0, r0
  404=>x"0612",	-- 0000011000010010  dec	r2, r2
  405=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  406=>x"FFF5",	-- 1111111111110101  liw	r5, paper_tilemap
  407=>x"17B0",	-- 0001011110110000  
  408=>x"D02C",	-- 1101000000101100  lw	r4, r5
  409=>x"042D",	-- 0000010000101101  inc	r5, r5
  410=>x"8960",	-- 1000100101100000  brieq	r4, PaperGameTileSkip
  411=>x"063F",	-- 0000011000111111  dec	r7, r7
  412=>x"D23D",	-- 1101001000111101  sw	r5, r7
  413=>x"FFF3",	-- 1111111111110011  liw	r3, paper_tilemap
  414=>x"17B0",	-- 0001011110110000  
  415=>x"0AEB",	-- 0000101011101011  sub	r3, r5, r3
  416=>x"6E20",	-- 0110111000100000  shr	r0, r4, 7
  417=>x"6219",	-- 0110001000011001  shr	r1, r3, 1
  418=>x"4809",	-- 0100100000001001  shl	r1, r1, 4
  419=>x"C19A",	-- 1100000110011010  li	r2, 51
  420=>x"0889",	-- 0000100010001001  add	r1, r1, r2
  421=>x"FFF2",	-- 1111111111110010  liw	r2, paper_pos + 1
  422=>x"179E",	-- 0001011110011110  
  423=>x"D012",	-- 1101000000010010  lw	r2, r2
  424=>x"6412",	-- 0110010000010010  shr	r2, r2, 2
  425=>x"C0FB",	-- 1100000011111011  li	r3, 31
  426=>x"20D2",	-- 0010000011010010  and	r2, r2, r3
  427=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  428=>x"4E24",	-- 0100111000100100  shl	r4, r4, 7
  429=>x"6E24",	-- 0110111000100100  shr	r4, r4, 7
  430=>x"C00B",	-- 1100000000001011  li	r3, 1
  431=>x"FB06",	-- 1111101100000110  bailne	r0, r6, put_tile
  432=>x"028D",	-- 0000001010001101  
  433=>x"81E0",	-- 1000000111100000  brieq	r4, PaperGameSegmentSkip
  435=>x"C013",	-- 1100000000010011  li	r3, 2
  436=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_tile
  437=>x"028D",	-- 0000001010001101  
  438=>x"0624",	-- 0000011000100100  dec	r4, r4
  439=>x"BF64",	-- 1011111101100100  brine	r4, PaperGameSegmentLoop
  440=>x"C003",	-- 1100000000000011  li	r3, 0
  441=>x"C144",	-- 1100000101000100  li	r4, 40
  442=>x"0B04",	-- 0000101100000100  sub	r4, r0, r4
  443=>x"FB66",	-- 1111101101100110  baillt	r4, r6, put_tile
  444=>x"028D",	-- 0000001010001101  
  445=>x"D03D",	-- 1101000000111101  lw	r5, r7
  446=>x"043F",	-- 0000010000111111  inc	r7, r7
  447=>x"FFF4",	-- 1111111111110100  liw r4, paper_tilemap + 24
  448=>x"17C8",	-- 0001011111001000  
  449=>x"0B2C",	-- 0000101100101100  sub	r4, r5, r4
  450=>x"B5A5",	-- 1011010110100101  brilt	r4, PaperGameTileLoop
  451=>x"FFF3",	-- 1111111111110011  liw	r3, paper_speed
  452=>x"17A0",	-- 0001011110100000  
  453=>x"D01B",	-- 1101000000011011  lw	r3, r3
  454=>x"CF84",	-- 1100111110000100  li	r4, 0x1F0
  455=>x"211C",	-- 0010000100011100  and	r4, r3, r4
  456=>x"FFF3",	-- 1111111111110011  liw	r3, paper_pos
  457=>x"179D",	-- 0001011110011101  
  458=>x"D018",	-- 1101000000011000  lw	r0, r3
  459=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  460=>x"FFF2",	-- 1111111111110010  liw	r2, paper_sprites
  461=>x"1720",	-- 0001011100100000  
  462=>x"0912",	-- 0000100100010010  add	r2, r2, r4
  463=>x"C161",	-- 1100000101100001  li	r1, 44
  464=>x"C083",	-- 1100000010000011  li	r3, 16
  465=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_16_masked
  466=>x"035D",	-- 0000001101011101  
  467=>x"902C",	-- 1001000000101100  brine	r5, PaperGameFail
  469=>x"C010",	-- 1100000000010000  li	r0, 2
  470=>x"C001",	-- 1100000000000001  li	r1, 0
  471=>x"8043",	-- 1000000001000011  bri	-, $+1
  472=>x"0609",	-- 0000011000001001  dec	r1, r1
  473=>x"BF8C",	-- 1011111110001100  brine	r1, $-2
  474=>x"0600",	-- 0000011000000000  dec	r0, r0
  475=>x"BEC4",	-- 1011111011000100  brine	r0, $-5
  476=>x"FFF2",	-- 1111111111110010  liw	r2, paper_pos
  477=>x"179D",	-- 0001011110011101  
  478=>x"FFF3",	-- 1111111111110011  liw	r3, paper_speed
  479=>x"17A0",	-- 0001011110100000  
  480=>x"D010",	-- 1101000000010000  lw	r0, r2
  481=>x"D019",	-- 1101000000011001  lw	r1, r3
  482=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  483=>x"8C05",	-- 1000110000000101  brilt	r0, PaperGameFail
  484=>x"FFF4",	-- 1111111111110100  liw	r4, 304*8
  485=>x"0980",	-- 0000100110000000  
  486=>x"0B04",	-- 0000101100000100  sub	r4, r0, r4
  487=>x"8B21",	-- 1000101100100001  brige	r4, PaperGameFail
  488=>x"D210",	-- 1101001000010000  sw	r0, r2
  489=>x"0412",	-- 0000010000010010  inc	r2, r2
  490=>x"041B",	-- 0000010000011011  inc	r3, r3
  491=>x"D010",	-- 1101000000010000  lw	r0, r2
  492=>x"D019",	-- 1101000000011001  lw	r1, r3
  493=>x"C7FC",	-- 1100011111111100  li	r4, 0xFF
  494=>x"6009",	-- 0110000000001001  shr	r1, r1, 0
  495=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  496=>x"2101",	-- 0010000100000001  and	r1, r0, r4
  497=>x"D211",	-- 1101001000010001  sw	r1, r2
  498=>x"2624",	-- 0010011000100100  not	r4, r4
  499=>x"2100",	-- 0010000100000000  and	r0, r0, r4
  500=>x"FB06",	-- 1111101100000110  bailne	r0, r6, PaperMapScroll
  501=>x"0235",	-- 0000001000110101  
  502=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  503=>x"16C0",	-- 0001011011000000  
  504=>x"D01B",	-- 1101000000011011  lw	r3, r3
  505=>x"F818",	-- 1111100000011000  baieq	r3, PaperGameRedraw
  506=>x"0144",	-- 0000000101000100  
  507=>x"F55C",	-- 1111010101011100  bspl	r4, r3, 5
  508=>x"8A24",	-- 1000101000100100  brine	r4, PaperGameQuit
  509=>x"F51C",	-- 1111010100011100  bspl	r4, r3, 4
  510=>x"89E4",	-- 1000100111100100  brine	r4, PaperGamePause
  511=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  512=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveUp
  513=>x"F49C",	-- 1111010010011100  bspl	r4, r3, 2
  514=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveDOWN
  515=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  516=>x"81A0",	-- 1000000110100000  brieq	r4, PaperNoMoveLEFT
  517=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  518=>x"17A0",	-- 0001011110100000  
  519=>x"D010",	-- 1101000000010000  lw	r0, r2
  520=>x"0600",	-- 0000011000000000  dec	r0, r0
  521=>x"D210",	-- 1101001000010000  sw	r0, r2
  522=>x"F4DC",	-- 1111010011011100  bspl	r4, r3, 3
  523=>x"81A0",	-- 1000000110100000  brieq	r4, PaperNoMoveRIGHT
  524=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  525=>x"17A0",	-- 0001011110100000  
  526=>x"D010",	-- 1101000000010000  lw	r0, r2
  527=>x"0400",	-- 0000010000000000  inc	r0, r0
  528=>x"D210",	-- 1101001000010000  sw	r0, r2
  529=>x"F8C0",	-- 1111100011000000  bai	-, PaperGameRedraw
  530=>x"0144",	-- 0000000101000100  
  531=>x"C000",	-- 1100000000000000  li	r0, 0
  532=>x"FFF2",	-- 1111111111110010  liw	r2, 240*20
  533=>x"12C0",	-- 0001001011000000  
  534=>x"D001",	-- 1101000000000001  lw	r1, r0
  535=>x"2609",	-- 0010011000001001  not	r1, r1
  536=>x"D201",	-- 1101001000000001  sw	r1, r0
  537=>x"0400",	-- 0000010000000000  inc	r0, r0
  538=>x"0612",	-- 0000011000010010  dec	r2, r2
  539=>x"BED4",	-- 1011111011010100  brine	r2, $-5
  540=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  541=>x"16C0",	-- 0001011011000000  
  542=>x"D01A",	-- 1101000000011010  lw	r2, r3
  543=>x"BFD4",	-- 1011111111010100  brine	r2, $-1
  544=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  545=>x"16C0",	-- 0001011011000000  
  546=>x"D01A",	-- 1101000000011010  lw	r2, r3
  547=>x"BFD0",	-- 1011111111010000  brieq	r2, $-1
  548=>x"FFFF",	-- 1111111111111111  reset
  549=>x"C080",	-- 1100000010000000  li	r0, 16
  550=>x"C0C1",	-- 1100000011000001  li	r1, 24
  551=>x"FFF2",	-- 1111111111110010  liw	r2, paper_pause
  552=>x"17C8",	-- 0001011111001000  
  553=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  554=>x"02BD",	-- 0000001010111101  
  555=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  556=>x"16C0",	-- 0001011011000000  
  557=>x"D01A",	-- 1101000000011010  lw	r2, r3
  558=>x"BFD4",	-- 1011111111010100  brine	r2, $-1
  559=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  560=>x"16C0",	-- 0001011011000000  
  561=>x"D01A",	-- 1101000000011010  lw	r2, r3
  562=>x"BFD0",	-- 1011111111010000  brieq	r2, $-1
  563=>x"F8C0",	-- 1111100011000000  bai	-, PaperGameRedraw
  564=>x"0144",	-- 0000000101000100  
  565=>x"FFF0",	-- 1111111111110000  liw	r0, paper_tilemap
  566=>x"17B0",	-- 0001011110110000  
  567=>x"C021",	-- 1100000000100001  li	r1, 4
  568=>x"0841",	-- 0000100001000001  add	r1, r0, r1
  569=>x"C0A2",	-- 1100000010100010  li	r2, 5*4
  570=>x"D00B",	-- 1101000000001011  lw	r3, r1
  571=>x"D203",	-- 1101001000000011  sw	r3, r0
  572=>x"0400",	-- 0000010000000000  inc	r0, r0
  573=>x"0409",	-- 0000010000001001  inc	r1, r1
  574=>x"0612",	-- 0000011000010010  dec	r2, r2
  575=>x"BED4",	-- 1011111011010100  brine	r2, PaperGameScrollLoop
  576=>x"063F",	-- 0000011000111111  dec	r7, r7
  577=>x"D23E",	-- 1101001000111110  sw	r6, r7
  578=>x"FAC6",	-- 1111101011000110  bail	-, r6, rand16
  579=>x"027B",	-- 0000001001111011  
  580=>x"C02A",	-- 1100000000101010  li	r2, 0x05
  581=>x"208B",	-- 0010000010001011  and	r3, r1, r2
  582=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  583=>x"208C",	-- 0010000010001100  and	r4, r1, r2
  584=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  585=>x"1F19",	-- 0001111100011001  mixll	r1, r3, r4
  586=>x"D201",	-- 1101001000000001  sw	r1, r0
  587=>x"0400",	-- 0000010000000000  inc	r0, r0
  588=>x"C03A",	-- 1100000000111010  li	r2, 0x07
  589=>x"091C",	-- 0000100100011100  add r4, r3, r4
  590=>x"208B",	-- 0010000010001011  and	r3, r1, r2
  591=>x"091C",	-- 0000100100011100  add r4, r3, r4
  592=>x"C01B",	-- 1100000000011011  li	r3, 3
  593=>x"08E4",	-- 0000100011100100  add	r4, r4, r3
  594=>x"6209",	-- 0110001000001001  shr	r1, r1, 1
  595=>x"208B",	-- 0010000010001011  and	r3, r1, r2
  596=>x"091B",	-- 0000100100011011  add r3, r3, r4
  597=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  598=>x"208C",	-- 0010000010001100  and	r4, r1, r2
  599=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  600=>x"1F19",	-- 0001111100011001  mixll	r1, r3, r4
  601=>x"D201",	-- 1101001000000001  sw	r1, r0
  602=>x"0400",	-- 0000010000000000  inc	r0, r0
  603=>x"C02A",	-- 1100000000101010  li	r2, 0x05
  604=>x"091C",	-- 0000100100011100  add r4, r3, r4
  605=>x"208B",	-- 0010000010001011  and	r3, r1, r2
  606=>x"091C",	-- 0000100100011100  add r4, r3, r4
  607=>x"C01B",	-- 1100000000011011  li	r3, 3
  608=>x"08E4",	-- 0000100011100100  add	r4, r4, r3
  609=>x"6209",	-- 0110001000001001  shr	r1, r1, 1
  610=>x"208B",	-- 0010000010001011  and	r3, r1, r2
  611=>x"091B",	-- 0000100100011011  add r3, r3, r4
  612=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  613=>x"208C",	-- 0010000010001100  and	r4, r1, r2
  614=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  615=>x"1F19",	-- 0001111100011001  mixll	r1, r3, r4
  616=>x"D201",	-- 1101001000000001  sw	r1, r0
  617=>x"0400",	-- 0000010000000000  inc	r0, r0
  618=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed + 1
  619=>x"17A1",	-- 0001011110100001  
  620=>x"D011",	-- 1101000000010001  lw	r1, r2
  621=>x"0409",	-- 0000010000001001  inc	r1, r1
  622=>x"D211",	-- 1101001000010001  sw	r1, r2
  623=>x"FFF2",	-- 1111111111110010  liw	r2, paper_score
  624=>x"16C9",	-- 0001011011001001  
  625=>x"D011",	-- 1101000000010001  lw	r1, r2
  626=>x"0409",	-- 0000010000001001  inc	r1, r1
  627=>x"D211",	-- 1101001000010001  sw	r1, r2
  628=>x"D03E",	-- 1101000000111110  lw	r6, r7
  629=>x"043F",	-- 0000010000111111  inc	r7, r7
  630=>x"E383",	-- 1110001110000011  ba	-, r6
  631=>x"FFF2",	-- 1111111111110010  liw	r2, rand_seed
  632=>x"16C8",	-- 0001011011001000  
  633=>x"D210",	-- 1101001000010000  sw	r0, r2
  634=>x"E383",	-- 1110001110000011  ba	-, r6
  635=>x"FFF2",	-- 1111111111110010  liw	r2, rand_seed
  636=>x"16C8",	-- 0001011011001000  
  637=>x"D013",	-- 1101000000010011  lw	r3, r2
  638=>x"C7EC",	-- 1100011111101100  li	r4, 253
  639=>x"1F19",	-- 0001111100011001  mixll	r1, r3, r4
  640=>x"18E4",	-- 0001100011100100  mixhh	r4, r4, r3
  641=>x"C002",	-- 1100000000000010  li	r2, 0
  642=>x"0AC9",	-- 0000101011001001  sub	r1, r1, r3
  643=>x"0EA4",	-- 0000111010100100  sbc	r4, r4, r2
  644=>x"0EC9",	-- 0000111011001001  sbc	r1, r1, r3
  645=>x"0EA4",	-- 0000111010100100  sbc	r4, r4, r2
  646=>x"1B13",	-- 0001101100010011  mixhl	r3, r2, r4
  647=>x"0EC9",	-- 0000111011001001  sbc	r1, r1, r3
  648=>x"0C89",	-- 0000110010001001  adc	r1, r1, r2
  649=>x"FFF2",	-- 1111111111110010  liw	r2, rand_seed
  650=>x"16C8",	-- 0001011011001000  
  651=>x"D211",	-- 1101001000010001  sw	r1, r2
  652=>x"E383",	-- 1110001110000011  ba	-, r6
  653=>x"063F",	-- 0000011000111111  dec	r7, r7
  654=>x"D238",	-- 1101001000111000  sw	r0, r7
  655=>x"063F",	-- 0000011000111111  dec	r7, r7
  656=>x"D239",	-- 1101001000111001  sw	r1, r7
  657=>x"063F",	-- 0000011000111111  dec	r7, r7
  658=>x"D23A",	-- 1101001000111010  sw	r2, r7
  659=>x"063F",	-- 0000011000111111  dec	r7, r7
  660=>x"D23B",	-- 1101001000111011  sw	r3, r7
  661=>x"063F",	-- 0000011000111111  dec	r7, r7
  662=>x"D23C",	-- 1101001000111100  sw	r4, r7
  663=>x"063F",	-- 0000011000111111  dec	r7, r7
  664=>x"D23D",	-- 1101001000111101  sw	r5, r7
  665=>x"063F",	-- 0000011000111111  dec	r7, r7
  666=>x"D23E",	-- 1101001000111110  sw	r6, r7
  667=>x"FFF2",	-- 1111111111110010  liw	r2, paper_tiles
  668=>x"1790",	-- 0001011110010000  
  669=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  670=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  671=>x"C043",	-- 1100000001000011  li	r3, 8
  672=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  673=>x"039F",	-- 0000001110011111  
  674=>x"D03E",	-- 1101000000111110  lw	r6, r7
  675=>x"043F",	-- 0000010000111111  inc	r7, r7
  676=>x"D03D",	-- 1101000000111101  lw	r5, r7
  677=>x"043F",	-- 0000010000111111  inc	r7, r7
  678=>x"D03C",	-- 1101000000111100  lw	r4, r7
  679=>x"043F",	-- 0000010000111111  inc	r7, r7
  680=>x"D03B",	-- 1101000000111011  lw	r3, r7
  681=>x"043F",	-- 0000010000111111  inc	r7, r7
  682=>x"D03A",	-- 1101000000111010  lw	r2, r7
  683=>x"043F",	-- 0000010000111111  inc	r7, r7
  684=>x"D039",	-- 1101000000111001  lw	r1, r7
  685=>x"043F",	-- 0000010000111111  inc	r7, r7
  686=>x"D038",	-- 1101000000111000  lw	r0, r7
  687=>x"043F",	-- 0000010000111111  inc	r7, r7
  688=>x"0400",	-- 0000010000000000  inc	r0, r0
  689=>x"E383",	-- 1110001110000011  ba	-, r6
  690=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  691=>x"C084",	-- 1100000010000100  li	r4, 16
  692=>x"0800",	-- 0000100000000000  add	r0, r0, r0
  693=>x"0C49",	-- 0000110001001001  adc	r1, r1, r1
  694=>x"0A8B",	-- 0000101010001011  sub	r3, r1, r2
  695=>x"80DD",	-- 1000000011011101  brilt	r3, div_16_16.skip
  696=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  697=>x"0400",	-- 0000010000000000  inc	r0, r0
  698=>x"0624",	-- 0000011000100100  dec	r4, r4
  699=>x"BE64",	-- 1011111001100100  brine	r4, div_16_16.loop
  700=>x"E383",	-- 1110001110000011  ba	-, r6
  701=>x"063F",	-- 0000011000111111  dec	r7, r7
  702=>x"D23E",	-- 1101001000111110  sw	r6, r7
  703=>x"D013",	-- 1101000000010011  lw	r3, r2
  704=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  705=>x"84D8",	-- 1000010011011000  brieq	r3, puts.end
  706=>x"063F",	-- 0000011000111111  dec	r7, r7
  707=>x"D23A",	-- 1101001000111010  sw	r2, r7
  708=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  709=>x"02D7",	-- 0000001011010111  
  710=>x"D03A",	-- 1101000000111010  lw	r2, r7
  711=>x"043F",	-- 0000010000111111  inc	r7, r7
  712=>x"D013",	-- 1101000000010011  lw	r3, r2
  713=>x"4E1B",	-- 0100111000011011  shl	r3, r3, 7
  714=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  715=>x"8258",	-- 1000001001011000  brieq	r3, puts.end
  716=>x"063F",	-- 0000011000111111  dec	r7, r7
  717=>x"D23A",	-- 1101001000111010  sw	r2, r7
  718=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  719=>x"02D7",	-- 0000001011010111  
  720=>x"D03A",	-- 1101000000111010  lw	r2, r7
  721=>x"043F",	-- 0000010000111111  inc	r7, r7
  722=>x"0412",	-- 0000010000010010  inc	r2, r2
  723=>x"BB03",	-- 1011101100000011  bri	-, puts.loop
  724=>x"D03E",	-- 1101000000111110  lw	r6, r7
  725=>x"043F",	-- 0000010000111111  inc	r7, r7
  726=>x"E383",	-- 1110001110000011  ba	-, r6
  727=>x"063F",	-- 0000011000111111  dec	r7, r7
  728=>x"D23E",	-- 1101001000111110  sw	r6, r7
  729=>x"063F",	-- 0000011000111111  dec	r7, r7
  730=>x"D238",	-- 1101001000111000  sw	r0, r7
  731=>x"063F",	-- 0000011000111111  dec	r7, r7
  732=>x"D239",	-- 1101001000111001  sw	r1, r7
  733=>x"FFF2",	-- 1111111111110010  liw	r2, font_map
  734=>x"12C0",	-- 0001001011000000  
  735=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  736=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  737=>x"C043",	-- 1100000001000011  li	r3, 8
  738=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  739=>x"039F",	-- 0000001110011111  
  740=>x"D039",	-- 1101000000111001  lw	r1, r7
  741=>x"043F",	-- 0000010000111111  inc	r7, r7
  742=>x"D038",	-- 1101000000111000  lw	r0, r7
  743=>x"043F",	-- 0000010000111111  inc	r7, r7
  744=>x"0400",	-- 0000010000000000  inc	r0, r0
  745=>x"D03E",	-- 1101000000111110  lw	r6, r7
  746=>x"043F",	-- 0000010000111111  inc	r7, r7
  747=>x"E383",	-- 1110001110000011  ba	-, r6
  748=>x"063F",	-- 0000011000111111  dec	r7, r7
  749=>x"D23E",	-- 1101001000111110  sw	r6, r7
  750=>x"FFF4",	-- 1111111111110100  liw	r4, 10000
  751=>x"2710",	-- 0010011100010000  
  752=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  753=>x"02FF",	-- 0000001011111111  
  754=>x"FFF4",	-- 1111111111110100  liw	r4, 1000
  755=>x"03E8",	-- 0000001111101000  
  756=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  757=>x"02FF",	-- 0000001011111111  
  758=>x"C324",	-- 1100001100100100  li	r4, 100
  759=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  760=>x"02FF",	-- 0000001011111111  
  761=>x"C054",	-- 1100000001010100  li	r4, 10
  762=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  763=>x"02FF",	-- 0000001011111111  
  764=>x"D03E",	-- 1101000000111110  lw	r6, r7
  765=>x"043F",	-- 0000010000111111  inc	r7, r7
  766=>x"C00C",	-- 1100000000001100  li	r4, 1
  767=>x"C17B",	-- 1100000101111011  li	r3, 0x2F
  768=>x"041B",	-- 0000010000011011  inc	r3, r3
  769=>x"0B12",	-- 0000101100010010  sub	r2, r2, r4
  770=>x"BF91",	-- 1011111110010001  brige	r2, printnum.loop
  771=>x"0912",	-- 0000100100010010  add	r2, r2, r4
  772=>x"063F",	-- 0000011000111111  dec	r7, r7
  773=>x"D23E",	-- 1101001000111110  sw	r6, r7
  774=>x"063F",	-- 0000011000111111  dec	r7, r7
  775=>x"D23A",	-- 1101001000111010  sw	r2, r7
  776=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  777=>x"02D7",	-- 0000001011010111  
  778=>x"D03A",	-- 1101000000111010  lw	r2, r7
  779=>x"043F",	-- 0000010000111111  inc	r7, r7
  780=>x"D03E",	-- 1101000000111110  lw	r6, r7
  781=>x"043F",	-- 0000010000111111  inc	r7, r7
  782=>x"E383",	-- 1110001110000011  ba	-, r6
  783=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  784=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  785=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  786=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  787=>x"C0A0",	-- 1100000010100000  li	r0, 20
  788=>x"0412",	-- 0000010000010010  inc	r2, r2
  789=>x"D011",	-- 1101000000010001  lw	r1, r2
  790=>x"E421",	-- 1110010000100001  exw	r1, r4
  791=>x"0412",	-- 0000010000010010  inc	r2, r2
  792=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  793=>x"061B",	-- 0000011000011011  dec	r3, r3
  794=>x"BE9C",	-- 1011111010011100  brine	r3, put_sprite_16_aligned.loop
  795=>x"C005",	-- 1100000000000101  li	r5, 0
  796=>x"E383",	-- 1110001110000011  ba	-, r6
  797=>x"C07D",	-- 1100000001111101  li	r5, 15
  798=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  799=>x"6600",	-- 0110011000000000  shr	r0, r0, 3
  800=>x"BBE8",	-- 1011101111101000  brieq	r5, put_sprite_16_aligned
  801=>x"062D",	-- 0000011000101101  dec	r5, r5
  802=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  803=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  804=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  805=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  806=>x"063F",	-- 0000011000111111  dec	r7, r7
  807=>x"D23B",	-- 1101001000111011  sw	r3, r7
  808=>x"0412",	-- 0000010000010010  inc	r2, r2
  809=>x"D011",	-- 1101000000010001  lw	r1, r2
  810=>x"CFF8",	-- 1100111111111000  li	r0, -1
  811=>x"3D40",	-- 0011110101000000  rsr	r0, r0, r5
  812=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  813=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  814=>x"D023",	-- 1101000000100011  lw	r3, r4
  815=>x"2600",	-- 0010011000000000  not	r0, r0
  816=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  817=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  818=>x"E421",	-- 1110010000100001  exw	r1, r4
  819=>x"0424",	-- 0000010000100100  inc	r4, r4
  820=>x"D011",	-- 1101000000010001  lw	r1, r2
  821=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  822=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  823=>x"D023",	-- 1101000000100011  lw	r3, r4
  824=>x"2600",	-- 0010011000000000  not	r0, r0
  825=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  826=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  827=>x"E421",	-- 1110010000100001  exw	r1, r4
  828=>x"0412",	-- 0000010000010010  inc	r2, r2
  829=>x"C098",	-- 1100000010011000  li	r0, 19
  830=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  831=>x"D03B",	-- 1101000000111011  lw	r3, r7
  832=>x"043F",	-- 0000010000111111  inc	r7, r7
  833=>x"061B",	-- 0000011000011011  dec	r3, r3
  834=>x"B91C",	-- 1011100100011100  brine	r3, put_sprite_16.loop
  835=>x"C005",	-- 1100000000000101  li	r5, 0
  836=>x"E383",	-- 1110001110000011  ba	-, r6
  837=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  838=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  839=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  840=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  841=>x"C005",	-- 1100000000000101  li	r5, 0
  842=>x"D020",	-- 1101000000100000  lw	r0, r4
  843=>x"D011",	-- 1101000000010001  lw	r1, r2
  844=>x"0412",	-- 0000010000010010  inc	r2, r2
  845=>x"2040",	-- 0010000001000000  and	r0, r0, r1
  846=>x"D011",	-- 1101000000010001  lw	r1, r2
  847=>x"2240",	-- 0010001001000000  or	r0, r0, r1
  848=>x"E420",	-- 1110010000100000  exw	r0, r4
  849=>x"0612",	-- 0000011000010010  dec	r2, r2
  850=>x"D011",	-- 1101000000010001  lw	r1, r2
  851=>x"2609",	-- 0010011000001001  not	r1, r1
  852=>x"0412",	-- 0000010000010010  inc	r2, r2
  853=>x"2040",	-- 0010000001000000  and	r0, r0, r1
  854=>x"222D",	-- 0010001000101101  or	r5, r5, r0
  855=>x"0412",	-- 0000010000010010  inc	r2, r2
  856=>x"C0A0",	-- 1100000010100000  li	r0, 20
  857=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  858=>x"061B",	-- 0000011000011011  dec	r3, r3
  859=>x"AE5C",	-- 1010111001011100  brine	r3, put_sprite_16_aligned.loop
  860=>x"E383",	-- 1110001110000011  ba	-, r6
  861=>x"C07D",	-- 1100000001111101  li	r5, 15
  862=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  863=>x"6600",	-- 0110011000000000  shr	r0, r0, 3
  864=>x"B968",	-- 1011100101101000  brieq	r5, put_sprite_16_masked_aligned
  865=>x"062D",	-- 0000011000101101  dec	r5, r5
  866=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  867=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  868=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  869=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  870=>x"063F",	-- 0000011000111111  dec	r7, r7
  871=>x"D23E",	-- 1101001000111110  sw	r6, r7
  872=>x"102E",	-- 0001000000101110  mova	r6, r5
  873=>x"C005",	-- 1100000000000101  li	r5, 0
  874=>x"063F",	-- 0000011000111111  dec	r7, r7
  875=>x"D23B",	-- 1101001000111011  sw	r3, r7
  876=>x"063F",	-- 0000011000111111  dec	r7, r7
  877=>x"D23D",	-- 1101001000111101  sw	r5, r7
  878=>x"D010",	-- 1101000000010000  lw	r0, r2
  879=>x"3980",	-- 0011100110000000  rrr	r0, r0, r6
  880=>x"0412",	-- 0000010000010010  inc	r2, r2
  881=>x"D011",	-- 1101000000010001  lw	r1, r2
  882=>x"3989",	-- 0011100110001001  rrr	r1, r1, r6
  883=>x"CFFD",	-- 1100111111111101  li	r5, -1
  884=>x"3DAD",	-- 0011110110101101  rsr	r5, r5, r6
  885=>x"2149",	-- 0010000101001001  and	r1, r1, r5
  886=>x"D023",	-- 1101000000100011  lw	r3, r4
  887=>x"262D",	-- 0010011000101101  not	r5, r5
  888=>x"222D",	-- 0010001000101101  or	r5, r5, r0
  889=>x"215B",	-- 0010000101011011  and	r3, r3, r5
  890=>x"225B",	-- 0010001001011011  or	r3, r3, r1
  891=>x"E423",	-- 1110010000100011  exw	r3, r4
  892=>x"262D",	-- 0010011000101101  not	r5, r5
  893=>x"215B",	-- 0010000101011011  and	r3, r3, r5
  894=>x"D03D",	-- 1101000000111101  lw	r5, r7
  895=>x"043F",	-- 0000010000111111  inc	r7, r7
  896=>x"22ED",	-- 0010001011101101  or	r5, r5, r3
  897=>x"0424",	-- 0000010000100100  inc	r4, r4
  898=>x"063F",	-- 0000011000111111  dec	r7, r7
  899=>x"D23D",	-- 1101001000111101  sw	r5, r7
  900=>x"D011",	-- 1101000000010001  lw	r1, r2
  901=>x"3989",	-- 0011100110001001  rrr	r1, r1, r6
  902=>x"CFFD",	-- 1100111111111101  li	r5, -1
  903=>x"3DAD",	-- 0011110110101101  rsr	r5, r5, r6
  904=>x"262D",	-- 0010011000101101  not	r5, r5
  905=>x"2149",	-- 0010000101001001  and	r1, r1, r5
  906=>x"D023",	-- 1101000000100011  lw	r3, r4
  907=>x"262D",	-- 0010011000101101  not	r5, r5
  908=>x"222D",	-- 0010001000101101  or	r5, r5, r0
  909=>x"215B",	-- 0010000101011011  and	r3, r3, r5
  910=>x"225B",	-- 0010001001011011  or	r3, r3, r1
  911=>x"E423",	-- 1110010000100011  exw	r3, r4
  912=>x"262D",	-- 0010011000101101  not	r5, r5
  913=>x"215B",	-- 0010000101011011  and	r3, r3, r5
  914=>x"D03D",	-- 1101000000111101  lw	r5, r7
  915=>x"043F",	-- 0000010000111111  inc	r7, r7
  916=>x"22ED",	-- 0010001011101101  or	r5, r5, r3
  917=>x"0412",	-- 0000010000010010  inc	r2, r2
  918=>x"C098",	-- 1100000010011000  li	r0, 19
  919=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  920=>x"D03B",	-- 1101000000111011  lw	r3, r7
  921=>x"043F",	-- 0000010000111111  inc	r7, r7
  922=>x"061B",	-- 0000011000011011  dec	r3, r3
  923=>x"B3DC",	-- 1011001111011100  brine	r3, put_sprite_16_masked.loop
  924=>x"D03E",	-- 1101000000111110  lw	r6, r7
  925=>x"043F",	-- 0000010000111111  inc	r7, r7
  926=>x"E383",	-- 1110001110000011  ba	-, r6
  927=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  928=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  929=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  930=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  931=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  932=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  933=>x"C0A5",	-- 1100000010100101  li	r5, 20
  934=>x"8404",	-- 1000010000000100  brine	r0, put_sprite_8_aligned.loop1
  935=>x"D010",	-- 1101000000010000  lw	r0, r2
  936=>x"D021",	-- 1101000000100001  lw	r1, r4
  937=>x"1A41",	-- 0001101001000001  mixhl	r1, r0, r1
  938=>x"D221",	-- 1101001000100001  sw	r1, r4
  939=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  940=>x"061B",	-- 0000011000011011  dec	r3, r3
  941=>x"E398",	-- 1110001110011000  baeq	r3, r6
  942=>x"D021",	-- 1101000000100001  lw	r1, r4
  943=>x"1E41",	-- 0001111001000001  mixll	r1, r0, r1
  944=>x"D221",	-- 1101001000100001  sw	r1, r4
  945=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  946=>x"0412",	-- 0000010000010010  inc	r2, r2
  947=>x"061B",	-- 0000011000011011  dec	r3, r3
  948=>x"E398",	-- 1110001110011000  baeq	r3, r6
  949=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop0
  950=>x"D010",	-- 1101000000010000  lw	r0, r2
  951=>x"D021",	-- 1101000000100001  lw	r1, r4
  952=>x"1809",	-- 0001100000001001  mixhh	r1, r1, r0
  953=>x"D221",	-- 1101001000100001  sw	r1, r4
  954=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  955=>x"061B",	-- 0000011000011011  dec	r3, r3
  956=>x"E398",	-- 1110001110011000  baeq	r3, r6
  957=>x"D021",	-- 1101000000100001  lw	r1, r4
  958=>x"1A09",	-- 0001101000001001  mixhl	r1, r1, r0
  959=>x"D221",	-- 1101001000100001  sw	r1, r4
  960=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  961=>x"0412",	-- 0000010000010010  inc	r2, r2
  962=>x"061B",	-- 0000011000011011  dec	r3, r3
  963=>x"E398",	-- 1110001110011000  baeq	r3, r6
  964=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop1
  965=>x"C03D",	-- 1100000000111101  li	r5, 7
  966=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  967=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  968=>x"B5E8",	-- 1011010111101000  brieq	r5, put_sprite_8_aligned
  969=>x"062D",	-- 0000011000101101  dec	r5, r5
  970=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  971=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  972=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  973=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  974=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  975=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  976=>x"8A04",	-- 1000101000000100  brine	r0, put_sprite_8.loop1
  977=>x"D010",	-- 1101000000010000  lw	r0, r2
  978=>x"063F",	-- 0000011000111111  dec	r7, r7
  979=>x"D23A",	-- 1101001000111010  sw	r2, r7
  980=>x"C802",	-- 1100100000000010  li	r2, 0x100
  981=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  982=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  983=>x"D021",	-- 1101000000100001  lw	r1, r4
  984=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  985=>x"2612",	-- 0010011000010010  not	r2, r2
  986=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  987=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  988=>x"D221",	-- 1101001000100001  sw	r1, r4
  989=>x"C0A1",	-- 1100000010100001  li	r1, 20
  990=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  991=>x"D03A",	-- 1101000000111010  lw	r2, r7
  992=>x"043F",	-- 0000010000111111  inc	r7, r7
  993=>x"061B",	-- 0000011000011011  dec	r3, r3
  994=>x"E398",	-- 1110001110011000  baeq	r3, r6
  995=>x"D010",	-- 1101000000010000  lw	r0, r2
  996=>x"063F",	-- 0000011000111111  dec	r7, r7
  997=>x"D23A",	-- 1101001000111010  sw	r2, r7
  998=>x"1E00",	-- 0001111000000000  mixll	r0, r0, r0
  999=>x"C802",	-- 1100100000000010  li	r2, 0x100
 1000=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
 1001=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
 1002=>x"D021",	-- 1101000000100001  lw	r1, r4
 1003=>x"2010",	-- 0010000000010000  and	r0, r2, r0
 1004=>x"2612",	-- 0010011000010010  not	r2, r2
 1005=>x"2089",	-- 0010000010001001  and	r1, r1, r2
 1006=>x"2209",	-- 0010001000001001  or	r1, r1, r0
 1007=>x"D221",	-- 1101001000100001  sw	r1, r4
 1008=>x"C0A1",	-- 1100000010100001  li	r1, 20
 1009=>x"0864",	-- 0000100001100100  add	r4, r4, r1
 1010=>x"D03A",	-- 1101000000111010  lw	r2, r7
 1011=>x"043F",	-- 0000010000111111  inc	r7, r7
 1012=>x"0412",	-- 0000010000010010  inc	r2, r2
 1013=>x"061B",	-- 0000011000011011  dec	r3, r3
 1014=>x"E398",	-- 1110001110011000  baeq	r3, r6
 1015=>x"B683",	-- 1011011010000011  bri	-, put_sprite_8.loop0
 1016=>x"D010",	-- 1101000000010000  lw	r0, r2
 1017=>x"063F",	-- 0000011000111111  dec	r7, r7
 1018=>x"D23A",	-- 1101001000111010  sw	r2, r7
 1019=>x"063F",	-- 0000011000111111  dec	r7, r7
 1020=>x"D23B",	-- 1101001000111011  sw	r3, r7
 1021=>x"C802",	-- 1100100000000010  li	r2, 0x100
 1022=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
 1023=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
 1024=>x"2080",	-- 0010000010000000  and	r0, r0, r2
 1025=>x"D021",	-- 1101000000100001  lw	r1, r4
 1026=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
 1027=>x"261B",	-- 0010011000011011  not	r3, r3
 1028=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
 1029=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
 1030=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
 1031=>x"D221",	-- 1101001000100001  sw	r1, r4
 1032=>x"0424",	-- 0000010000100100  inc	r4, r4
 1033=>x"D021",	-- 1101000000100001  lw	r1, r4
 1034=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
 1035=>x"261B",	-- 0010011000011011  not	r3, r3
 1036=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
 1037=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
 1038=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
 1039=>x"D221",	-- 1101001000100001  sw	r1, r4
 1040=>x"C099",	-- 1100000010011001  li	r1, 19
 1041=>x"0864",	-- 0000100001100100  add	r4, r4, r1
 1042=>x"D03B",	-- 1101000000111011  lw	r3, r7
 1043=>x"043F",	-- 0000010000111111  inc	r7, r7
 1044=>x"D03A",	-- 1101000000111010  lw	r2, r7
 1045=>x"043F",	-- 0000010000111111  inc	r7, r7
 1046=>x"061B",	-- 0000011000011011  dec	r3, r3
 1047=>x"E398",	-- 1110001110011000  baeq	r3, r6
 1048=>x"D010",	-- 1101000000010000  lw	r0, r2
 1049=>x"4E00",	-- 0100111000000000  shl	r0, r0, 7
 1050=>x"063F",	-- 0000011000111111  dec	r7, r7
 1051=>x"D23A",	-- 1101001000111010  sw	r2, r7
 1052=>x"063F",	-- 0000011000111111  dec	r7, r7
 1053=>x"D23B",	-- 1101001000111011  sw	r3, r7
 1054=>x"C802",	-- 1100100000000010  li	r2, 0x100
 1055=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
 1056=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
 1057=>x"2080",	-- 0010000010000000  and	r0, r0, r2
 1058=>x"D021",	-- 1101000000100001  lw	r1, r4
 1059=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
 1060=>x"261B",	-- 0010011000011011  not	r3, r3
 1061=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
 1062=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
 1063=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
 1064=>x"D221",	-- 1101001000100001  sw	r1, r4
 1065=>x"0424",	-- 0000010000100100  inc	r4, r4
 1066=>x"D021",	-- 1101000000100001  lw	r1, r4
 1067=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
 1068=>x"261B",	-- 0010011000011011  not	r3, r3
 1069=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
 1070=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
 1071=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
 1072=>x"D221",	-- 1101001000100001  sw	r1, r4
 1073=>x"C099",	-- 1100000010011001  li	r1, 19
 1074=>x"0864",	-- 0000100001100100  add	r4, r4, r1
 1075=>x"D03B",	-- 1101000000111011  lw	r3, r7
 1076=>x"043F",	-- 0000010000111111  inc	r7, r7
 1077=>x"D03A",	-- 1101000000111010  lw	r2, r7
 1078=>x"043F",	-- 0000010000111111  inc	r7, r7
 1079=>x"0412",	-- 0000010000010010  inc	r2, r2
 1080=>x"061B",	-- 0000011000011011  dec	r3, r3
 1081=>x"E398",	-- 1110001110011000  baeq	r3, r6
 1082=>x"AF83",	-- 1010111110000011  bri	-, put_sprite_8.loop1
    others => x"0000"
    );
begin
  process(CLK)
  begin
    if (CLK'event AND CLK='1') then
      D <= m(to_integer(unsigned(AD)));
    end if;
  end process;
end Behavioral;
