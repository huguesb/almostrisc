----------------------------------------------------------------------------------
--
-- File retrieved, on 07/02/2010, from :
-- http://sebastien-viardot.imag.fr/Enseignements/Archi1A2s/sources/ROMPROG.vhd
--
-- Slightly altered to get rid of vendor-specific packages and adjust formatting
-- Now auto-filled by asrom script
--
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROMPROG is
  Port ( AD : in  STD_LOGIC_VECTOR (12 downto 0);
         D : out  STD_LOGIC_VECTOR (15 downto 0);
         CLK : in STD_LOGIC);
end ROMPROG;

architecture Behavioral of ROMPROG is
  constant low_address: natural := 0;
  constant high_address: natural := 8192;
  subtype octet is std_logic_vector( 15 downto 0 );
  type zone_memoire is
    array (natural range low_address to high_address-1) of octet;
  constant m: zone_memoire:= (
    0=>x"FFF7",	-- 1111111111110111  liw	r7, IRQ_mask
    1=>x"2000",	-- 0010000000000000  
    2=>x"F8C0",	-- 1111100011000000  bai	-, os_init
    3=>x"0100",	-- 0000000100000000  
   16=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_ack
   17=>x"2002",	-- 0010000000000010  
   18=>x"D001",	-- 1101000000000001  lw	r1, r0
   19=>x"F54A",	-- 1111010101001010  bspl	r2, r1, 5
   20=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_error
   21=>x"0050",	-- 0000000001010000  
   22=>x"F4CA",	-- 1111010011001010  bspl	r2, r1, 3
   23=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_kbd
   24=>x"0060",	-- 0000000001100000  
   25=>x"F40A",	-- 1111010000001010  bspl	r2, r1, 0
   26=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_tmr
   27=>x"0040",	-- 0000000001000000  
   28=>x"D201",	-- 1101001000000001  sw	r1, r0
   29=>x"FFFE",	-- 1111111111111110  reti
   64=>x"263F",	-- 0010011000111111  not r7, r7
   65=>x"D7C0",	-- 1101011111000000  out	r7
   66=>x"E383",	-- 1110001110000011  ba	-, r6
   80=>x"25FF",	-- 0010010111111111  xor	r7, r7, r7
   81=>x"D7C0",	-- 1101011111000000  out	r7
   82=>x"E383",	-- 1110001110000011  ba	-, r6
   96=>x"FFF2",	-- 1111111111110010  liw	r2, PS2_rx
   97=>x"2004",	-- 0010000000000100  
   98=>x"D012",	-- 1101000000010010  lw	r2, r2
   99=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map + 8
  100=>x"1808",	-- 0001100000001000  
  101=>x"D01B",	-- 1101000000011011  lw	r3, r3
  102=>x"1EBF",	-- 0001111010111111  mixll	r7, r7, r2
  103=>x"C784",	-- 1100011110000100  li	r4, 0xF0
  104=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  105=>x"8B20",	-- 1000101100100000  brieq	r4, int_kbd.release
  106=>x"C704",	-- 1100011100000100  li	r4, 0xE0
  107=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  108=>x"88E0",	-- 1000100011100000  brieq	r4, int_kbd.extended
  109=>x"FFF5",	-- 1111111111110101  liw	r5, paper_keys - 1
  110=>x"16BF",	-- 0001011010111111  
  111=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  112=>x"80E0",	-- 1000000011100000  brieq	r4, $+3
  113=>x"FFF5",	-- 1111111111110101  liw	r5, paper_keys + 11 - 1
  114=>x"16CA",	-- 0001011011001010  
  115=>x"042D",	-- 0000010000101101  inc	r5, r5
  116=>x"D02C",	-- 1101000000101100  lw	r4, r5
  117=>x"8560",	-- 1000010101100000  brieq	r4, scan_code_mismatch
  118=>x"6E24",	-- 0110111000100100  shr	r4, r4, 7
  119=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  120=>x"BEE4",	-- 1011111011100100  brine	r4, scan_code_loop
  121=>x"D02A",	-- 1101000000101010  lw	r2, r5
  122=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  123=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  124=>x"741B",	-- 0111010000011011  shr	r3, r3, 10
  125=>x"C00D",	-- 1100000000001101  li	r5, 1
  126=>x"0612",	-- 0000011000010010  dec	r2, r2
  127=>x"3AAA",	-- 0011101010101010  rrl	r2, r5, r2
  128=>x"FFF5",	-- 1111111111110101  liw	r5, key_press_map
  129=>x"1800",	-- 0001100000000000  
  130=>x"08ED",	-- 0000100011101101  add	r5, r5, r3
  131=>x"D02B",	-- 1101000000101011  lw	r3, r5
  132=>x"80E4",	-- 1000000011100100  brine	r4, scan_code_release
  133=>x"229B",	-- 0010001010011011  or	r3, r3, r2
  134=>x"80C3",	-- 1000000011000011  bri	-, scan_code_notify
  135=>x"2612",	-- 0010011000010010  not	r2, r2
  136=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  137=>x"D22B",	-- 1101001000101011  sw	r3, r5
  138=>x"C003",	-- 1100000000000011  li	r3, 0
  139=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  140=>x"1808",	-- 0001100000001000  
  141=>x"D223",	-- 1101001000100011  sw	r3, r4
  142=>x"E383",	-- 1110001110000011  ba	-, r6
  143=>x"C014",	-- 1100000000010100  li	r4, 2
  144=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  145=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  146=>x"1808",	-- 0001100000001000  
  147=>x"D223",	-- 1101001000100011  sw	r3, r4
  148=>x"E383",	-- 1110001110000011  ba	-, r6
  149=>x"C00C",	-- 1100000000001100  li	r4, 1
  150=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  151=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  152=>x"1808",	-- 0001100000001000  
  153=>x"D223",	-- 1101001000100011  sw	r3, r4
  154=>x"E383",	-- 1110001110000011  ba	-, r6
  256=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_mask
  257=>x"2000",	-- 0010000000000000  
  258=>x"C0C9",	-- 1100000011001001  li	r1, 0x19
  259=>x"D201",	-- 1101001000000001  sw	r1, r0
  260=>x"0400",	-- 0000010000000000  inc	r0, r0
  261=>x"CFF9",	-- 1100111111111001  li	r1, -1
  262=>x"D201",	-- 1101001000000001  sw	r1, r0
  263=>x"C03A",	-- 1100000000111010  li	r2, 7
  264=>x"0880",	-- 0000100010000000  add	r0, r0, r2
  265=>x"C0EA",	-- 1100000011101010  li	r2, 0x1D
  266=>x"D202",	-- 1101001000000010  sw	r2, r0
  267=>x"0400",	-- 0000010000000000  inc	r0, r0
  268=>x"C07A",	-- 1100000001111010  li	r2, 15
  269=>x"D202",	-- 1101001000000010  sw	r2, r0
  270=>x"FFF0",	-- 1111111111110000  liw	r0, key_press_map
  271=>x"1800",	-- 0001100000000000  
  272=>x"C001",	-- 1100000000000001  li	r1, 0
  273=>x"C042",	-- 1100000001000010  li	r2, 8
  274=>x"D201",	-- 1101001000000001  sw	r1, r0
  275=>x"0400",	-- 0000010000000000  inc	r0, r0
  276=>x"0612",	-- 0000011000010010  dec	r2, r2
  277=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  278=>x"C0F3",	-- 1100000011110011  li	r3, 30
  279=>x"CFFA",	-- 1100111111111010  li	r2, -1
  280=>x"D21A",	-- 1101001000011010  sw	r2, r3
  281=>x"8083",	-- 1000000010000011  bri	-, PaperGameStart
  282=>x"8003",	-- 1000000000000011  bri	-, PaperMenuLoop
  283=>x"FFF0",	-- 1111111111110000  liw	r0, paper_dir
  284=>x"173C",	-- 0001011100111100  
  285=>x"C001",	-- 1100000000000001  li	r1, 0
  286=>x"D201",	-- 1101001000000001  sw	r1, r0
  287=>x"0400",	-- 0000010000000000  inc	r0, r0
  288=>x"FFF1",	-- 1111111111110001  liw	r1, 152 * 8
  289=>x"04C0",	-- 0000010011000000  
  290=>x"D201",	-- 1101001000000001  sw	r1, r0
  291=>x"0400",	-- 0000010000000000  inc	r0, r0
  292=>x"C001",	-- 1100000000000001  li	r1, 0
  293=>x"D201",	-- 1101001000000001  sw	r1, r0
  294=>x"0400",	-- 0000010000000000  inc	r0, r0
  295=>x"FFF1",	-- 1111111111110001  liw	r1, 128 * 8
  296=>x"0400",	-- 0000010000000000  
  297=>x"D201",	-- 1101001000000001  sw	r1, r0
  298=>x"0400",	-- 0000010000000000  inc	r0, r0
  299=>x"C001",	-- 1100000000000001  li	r1, 0
  300=>x"D201",	-- 1101001000000001  sw	r1, r0
  301=>x"0400",	-- 0000010000000000  inc	r0, r0
  302=>x"C029",	-- 1100000000101001  li	r1, 5
  303=>x"D201",	-- 1101001000000001  sw	r1, r0
  304=>x"0400",	-- 0000010000000000  inc	r0, r0
  305=>x"C011",	-- 1100000000010001  li	r1, 2
  306=>x"D201",	-- 1101001000000001  sw	r1, r0
  307=>x"0400",	-- 0000010000000000  inc	r0, r0
  308=>x"C000",	-- 1100000000000000  li	r0, 0
  309=>x"CFF9",	-- 1100111111111001  li	r1, -1
  310=>x"C0A2",	-- 1100000010100010  li	r2, 20
  311=>x"D201",	-- 1101001000000001  sw	r1, r0
  312=>x"0400",	-- 0000010000000000  inc	r0, r0
  313=>x"0612",	-- 0000011000010010  dec	r2, r2
  314=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  315=>x"C001",	-- 1100000000000001  li	r1, 0
  316=>x"FFF2",	-- 1111111111110010  liw	r2, 18*20
  317=>x"0168",	-- 0000000101101000  
  318=>x"D201",	-- 1101001000000001  sw	r1, r0
  319=>x"0400",	-- 0000010000000000  inc	r0, r0
  320=>x"0612",	-- 0000011000010010  dec	r2, r2
  321=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  322=>x"CFF9",	-- 1100111111111001  li	r1, -1
  323=>x"C0A2",	-- 1100000010100010  li	r2, 20
  324=>x"D201",	-- 1101001000000001  sw	r1, r0
  325=>x"0400",	-- 0000010000000000  inc	r0, r0
  326=>x"0612",	-- 0000011000010010  dec	r2, r2
  327=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  328=>x"C020",	-- 1100000000100000  li	r0, 4
  329=>x"C029",	-- 1100000000101001  li	r1, 5
  330=>x"FFF2",	-- 1111111111110010  liw	r2, paper_title
  331=>x"1744",	-- 0001011101000100  
  332=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  333=>x"0251",	-- 0000001001010001  
  334=>x"C778",	-- 1100011101111000  li	r0, 239
  335=>x"C009",	-- 1100000000001001  li	r1, 1
  336=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud
  337=>x"1720",	-- 0001011100100000  
  338=>x"C043",	-- 1100000001000011  li	r3, 8
  339=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  340=>x"02FB",	-- 0000001011111011  
  341=>x"C0F8",	-- 1100000011111000  li	r0, 31
  342=>x"C009",	-- 1100000000001001  li	r1, 1
  343=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed + 1
  344=>x"1741",	-- 0001011101000001  
  345=>x"D012",	-- 1101000000010010  lw	r2, r2
  346=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum
  347=>x"0280",	-- 0000001010000000  
  348=>x"C120",	-- 1100000100100000  li	r0, 36
  349=>x"C009",	-- 1100000000001001  li	r1, 1
  350=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  351=>x"174A",	-- 0001011101001010  
  352=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  353=>x"0251",	-- 0000001001010001  
  354=>x"C778",	-- 1100011101111000  li	r0, 239
  355=>x"C051",	-- 1100000001010001  li	r1, 10
  356=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud + 4
  357=>x"1724",	-- 0001011100100100  
  358=>x"C043",	-- 1100000001000011  li	r3, 8
  359=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  360=>x"02FB",	-- 0000001011111011  
  361=>x"C0F8",	-- 1100000011111000  li	r0, 31
  362=>x"C051",	-- 1100000001010001  li	r1, 10
  363=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed + 2
  364=>x"1742",	-- 0001011101000010  
  365=>x"D012",	-- 1101000000010010  lw	r2, r2
  366=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum
  367=>x"0280",	-- 0000001010000000  
  368=>x"C120",	-- 1100000100100000  li	r0, 36
  369=>x"C051",	-- 1100000001010001  li	r1, 10
  370=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  371=>x"174A",	-- 0001011101001010  
  372=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  373=>x"0251",	-- 0000001001010001  
  374=>x"FFF0",	-- 1111111111110000  liw	r0, 20*20
  375=>x"0190",	-- 0000000110010000  
  376=>x"C001",	-- 1100000000000001  li	r1, 0
  377=>x"FFF2",	-- 1111111111110010  liw	r2, 220*20
  378=>x"1130",	-- 0001000100110000  
  379=>x"D201",	-- 1101001000000001  sw	r1, r0
  380=>x"0400",	-- 0000010000000000  inc	r0, r0
  381=>x"0612",	-- 0000011000010010  dec	r2, r2
  382=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  383=>x"FFF5",	-- 1111111111110101  liw	r5, paper_tilemap
  384=>x"1780",	-- 0001011110000000  
  385=>x"D02C",	-- 1101000000101100  lw	r4, r5
  386=>x"042D",	-- 0000010000101101  inc	r5, r5
  387=>x"88E0",	-- 1000100011100000  brieq	r4, PaperGameTileSkip
  388=>x"063F",	-- 0000011000111111  dec	r7, r7
  389=>x"D23D",	-- 1101001000111101  sw	r5, r7
  390=>x"FFF3",	-- 1111111111110011  liw	r3, paper_tilemap
  391=>x"1780",	-- 0001011110000000  
  392=>x"0AEB",	-- 0000101011101011  sub	r3, r5, r3
  393=>x"6E20",	-- 0110111000100000  shr	r0, r4, 7
  394=>x"6219",	-- 0110001000011001  shr	r1, r3, 1
  395=>x"4409",	-- 0100010000001001  shl	r1, r1, 2
  396=>x"C0C2",	-- 1100000011000010  li	r2, 24
  397=>x"0889",	-- 0000100010001001  add	r1, r1, r2
  398=>x"FFF2",	-- 1111111111110010  liw	r2, paper_pos + 1
  399=>x"173E",	-- 0001011100111110  
  400=>x"D012",	-- 1101000000010010  lw	r2, r2
  401=>x"6412",	-- 0110010000010010  shr	r2, r2, 2
  402=>x"C03B",	-- 1100000000111011  li	r3, 7
  403=>x"20D2",	-- 0010000011010010  and	r2, r2, r3
  404=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  405=>x"4E24",	-- 0100111000100100  shl	r4, r4, 7
  406=>x"6E24",	-- 0110111000100100  shr	r4, r4, 7
  407=>x"C00B",	-- 1100000000001011  li	r3, 1
  408=>x"FB06",	-- 1111101100000110  bailne	r0, r6, put_tile
  409=>x"01FD",	-- 0000000111111101  
  410=>x"C013",	-- 1100000000010011  li	r3, 2
  411=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_tile
  412=>x"01FD",	-- 0000000111111101  
  413=>x"0624",	-- 0000011000100100  dec	r4, r4
  414=>x"BF64",	-- 1011111101100100  brine	r4, PaperGameSegmentLoop
  415=>x"C003",	-- 1100000000000011  li	r3, 0
  416=>x"C144",	-- 1100000101000100  li	r4, 40
  417=>x"0B04",	-- 0000101100000100  sub	r4, r0, r4
  418=>x"FB66",	-- 1111101101100110  baillt	r4, r6, put_tile
  419=>x"01FD",	-- 0000000111111101  
  420=>x"D03D",	-- 1101000000111101  lw	r5, r7
  421=>x"043F",	-- 0000010000111111  inc	r7, r7
  422=>x"FFF4",	-- 1111111111110100  liw r4, paper_tilemap + 125
  423=>x"17FD",	-- 0001011111111101  
  424=>x"0B2C",	-- 0000101100101100  sub	r4, r5, r4
  425=>x"B625",	-- 1011011000100101  brilt	r4, PaperGameTileLoop
  426=>x"FFF3",	-- 1111111111110011  liw	r3, paper_speed
  427=>x"1740",	-- 0001011101000000  
  428=>x"D01C",	-- 1101000000011100  lw	r4, r3
  429=>x"F7E5",	-- 1111011111100101  bspl	r5, r4, 15
  430=>x"2564",	-- 0010010101100100  xor	r4, r4, r5
  431=>x"6424",	-- 0110010000100100  shr	r4, r4, 2
  432=>x"2564",	-- 0010010101100100  xor	r4, r4, r5
  433=>x"FFF3",	-- 1111111111110011  liw	r3, paper_pos
  434=>x"173D",	-- 0001011100111101  
  435=>x"D018",	-- 1101000000011000  lw	r0, r3
  436=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  437=>x"FFF2",	-- 1111111111110010  liw	r2, paper_sprites
  438=>x"16F0",	-- 0001011011110000  
  439=>x"4624",	-- 0100011000100100  shl	r4, r4, 3
  440=>x"0912",	-- 0000100100010010  add	r2, r2, r4
  441=>x"C161",	-- 1100000101100001  li	r1, 44
  442=>x"C083",	-- 1100000010000011  li	r3, 16
  443=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_16
  444=>x"02AF",	-- 0000001010101111  
  445=>x"C028",	-- 1100000000101000  li	r0, 5
  446=>x"C001",	-- 1100000000000001  li	r1, 0
  447=>x"8043",	-- 1000000001000011  bri	-, $+1
  448=>x"8043",	-- 1000000001000011  bri	-, $+1
  449=>x"0609",	-- 0000011000001001  dec	r1, r1
  450=>x"BF4C",	-- 1011111101001100  brine	r1, $-3
  451=>x"0600",	-- 0000011000000000  dec	r0, r0
  452=>x"BE84",	-- 1011111010000100  brine	r0, $-6
  453=>x"FFF2",	-- 1111111111110010  liw	r2, paper_pos
  454=>x"173D",	-- 0001011100111101  
  455=>x"FFF3",	-- 1111111111110011  liw	r3, paper_speed
  456=>x"1740",	-- 0001011101000000  
  457=>x"D010",	-- 1101000000010000  lw	r0, r2
  458=>x"D019",	-- 1101000000011001  lw	r1, r3
  459=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  460=>x"D210",	-- 1101001000010000  sw	r0, r2
  461=>x"0412",	-- 0000010000010010  inc	r2, r2
  462=>x"041B",	-- 0000010000011011  inc	r3, r3
  463=>x"D010",	-- 1101000000010000  lw	r0, r2
  464=>x"D019",	-- 1101000000011001  lw	r1, r3
  465=>x"C1FC",	-- 1100000111111100  li	r4, 0x3F
  466=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  467=>x"2101",	-- 0010000100000001  and	r1, r0, r4
  468=>x"2624",	-- 0010011000100100  not	r4, r4
  469=>x"2100",	-- 0010000100000000  and	r0, r0, r4
  470=>x"D211",	-- 1101001000010001  sw	r1, r2
  471=>x"8300",	-- 1000001100000000  brieq	r0, PaperGameSkipScroll
  472=>x"FFF0",	-- 1111111111110000  liw	r0, paper_tilemap
  473=>x"1780",	-- 0001011110000000  
  474=>x"C021",	-- 1100000000100001  li	r1, 4
  475=>x"0841",	-- 0000100001000001  add	r1, r0, r1
  476=>x"C302",	-- 1100001100000010  li	r2, 24*4
  477=>x"D00B",	-- 1101000000001011  lw	r3, r1
  478=>x"D203",	-- 1101001000000011  sw	r3, r0
  479=>x"0400",	-- 0000010000000000  inc	r0, r0
  480=>x"0409",	-- 0000010000001001  inc	r1, r1
  481=>x"0612",	-- 0000011000010010  dec	r2, r2
  482=>x"BED4",	-- 1011111011010100  brine	r2, PaperGameScrollLoop
  483=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  484=>x"1800",	-- 0001100000000000  
  485=>x"D01B",	-- 1101000000011011  lw	r3, r3
  486=>x"A418",	-- 1010010000011000  brieq	r3, PaperGameRedrawContent
  487=>x"F7DC",	-- 1111011111011100  bspl	r4, r3, 15
  488=>x"8524",	-- 1000010100100100  brine	r4, PaperGameQuit
  489=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  490=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveUp
  491=>x"F49C",	-- 1111010010011100  bspl	r4, r3, 2
  492=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveDOWN
  493=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  494=>x"81A0",	-- 1000000110100000  brieq	r4, PaperNoMoveLEFT
  495=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  496=>x"1740",	-- 0001011101000000  
  497=>x"D010",	-- 1101000000010000  lw	r0, r2
  498=>x"0600",	-- 0000011000000000  dec	r0, r0
  499=>x"D210",	-- 1101001000010000  sw	r0, r2
  500=>x"F4DC",	-- 1111010011011100  bspl	r4, r3, 3
  501=>x"81A0",	-- 1000000110100000  brieq	r4, PaperNoMoveRIGHT
  502=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  503=>x"1740",	-- 0001011101000000  
  504=>x"D010",	-- 1101000000010000  lw	r0, r2
  505=>x"0400",	-- 0000010000000000  inc	r0, r0
  506=>x"D210",	-- 1101001000010000  sw	r0, r2
  507=>x"9EC3",	-- 1001111011000011  bri	-, PaperGameRedrawContent
  508=>x"FFFF",	-- 1111111111111111  reset
  509=>x"063F",	-- 0000011000111111  dec	r7, r7
  510=>x"D238",	-- 1101001000111000  sw	r0, r7
  511=>x"063F",	-- 0000011000111111  dec	r7, r7
  512=>x"D239",	-- 1101001000111001  sw	r1, r7
  513=>x"063F",	-- 0000011000111111  dec	r7, r7
  514=>x"D23A",	-- 1101001000111010  sw	r2, r7
  515=>x"063F",	-- 0000011000111111  dec	r7, r7
  516=>x"D23B",	-- 1101001000111011  sw	r3, r7
  517=>x"063F",	-- 0000011000111111  dec	r7, r7
  518=>x"D23C",	-- 1101001000111100  sw	r4, r7
  519=>x"063F",	-- 0000011000111111  dec	r7, r7
  520=>x"D23D",	-- 1101001000111101  sw	r5, r7
  521=>x"063F",	-- 0000011000111111  dec	r7, r7
  522=>x"D23E",	-- 1101001000111110  sw	r6, r7
  523=>x"FFF2",	-- 1111111111110010  liw	r2, paper_tiles
  524=>x"1730",	-- 0001011100110000  
  525=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  526=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  527=>x"C043",	-- 1100000001000011  li	r3, 8
  528=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  529=>x"02D5",	-- 0000001011010101  
  530=>x"D03E",	-- 1101000000111110  lw	r6, r7
  531=>x"043F",	-- 0000010000111111  inc	r7, r7
  532=>x"D03D",	-- 1101000000111101  lw	r5, r7
  533=>x"043F",	-- 0000010000111111  inc	r7, r7
  534=>x"D03C",	-- 1101000000111100  lw	r4, r7
  535=>x"043F",	-- 0000010000111111  inc	r7, r7
  536=>x"D03B",	-- 1101000000111011  lw	r3, r7
  537=>x"043F",	-- 0000010000111111  inc	r7, r7
  538=>x"D03A",	-- 1101000000111010  lw	r2, r7
  539=>x"043F",	-- 0000010000111111  inc	r7, r7
  540=>x"D039",	-- 1101000000111001  lw	r1, r7
  541=>x"043F",	-- 0000010000111111  inc	r7, r7
  542=>x"D038",	-- 1101000000111000  lw	r0, r7
  543=>x"043F",	-- 0000010000111111  inc	r7, r7
  544=>x"0400",	-- 0000010000000000  inc	r0, r0
  545=>x"E383",	-- 1110001110000011  ba	-, r6
  546=>x"C750",	-- 1100011101010000  li	r0, 234
  547=>x"C1C2",	-- 1100000111000010  li	r2, 56
  548=>x"FAC6",	-- 1111101011000110  bail	-, r6, div_16_16
  549=>x"023A",	-- 0000001000111010  
  550=>x"C448",	-- 1100010001001000  li	r0, 137
  551=>x"C472",	-- 1100010001110010  li	r2, 142
  552=>x"FAC6",	-- 1111101011000110  bail	-, r6, mult_16_16
  553=>x"022E",	-- 0000001000101110  
  554=>x"C03A",	-- 1100000000111010  li r2, 7
  555=>x"FAC6",	-- 1111101011000110  bail	-, r6, fact_16
  556=>x"0245",	-- 0000001001000101  
  557=>x"FFFF",	-- 1111111111111111  reset
  558=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  559=>x"2524",	-- 0010010100100100  xor	r4, r4, r4
  560=>x"C085",	-- 1100000010000101  li	r5, 16
  561=>x"0849",	-- 0000100001001001  add	r1, r1, r1
  562=>x"0C00",	-- 0000110000000000  adc	r0, r0, r0
  563=>x"0EDB",	-- 0000111011011011  sbc	r3, r3, r3
  564=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  565=>x"08C9",	-- 0000100011001001  add	r1, r1, r3
  566=>x"0D00",	-- 0000110100000000  adc	r0, r0, r4
  567=>x"062D",	-- 0000011000101101  dec	r5, r5
  568=>x"BE6C",	-- 1011111001101100  brine	r5, mult_16_16.loop
  569=>x"E383",	-- 1110001110000011  ba	-, r6
  570=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  571=>x"C084",	-- 1100000010000100  li	r4, 16
  572=>x"0800",	-- 0000100000000000  add	r0, r0, r0
  573=>x"0C49",	-- 0000110001001001  adc	r1, r1, r1
  574=>x"0A8B",	-- 0000101010001011  sub	r3, r1, r2
  575=>x"80DD",	-- 1000000011011101  brilt	r3, div_16_16.skip
  576=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  577=>x"0400",	-- 0000010000000000  inc	r0, r0
  578=>x"0624",	-- 0000011000100100  dec	r4, r4
  579=>x"BE64",	-- 1011111001100100  brine	r4, div_16_16.loop
  580=>x"E383",	-- 1110001110000011  ba	-, r6
  581=>x"2400",	-- 0010010000000000  xor	r0, r0, r0
  582=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  583=>x"8250",	-- 1000001001010000  brieq	r2, fact_16.end
  584=>x"0409",	-- 0000010000001001  inc	r1, r1
  585=>x"1008",	-- 0001000000001000  mova	r0, r1
  586=>x"FAC6",	-- 1111101011000110  bail	-, r6, mult_16_16
  587=>x"022E",	-- 0000001000101110  
  588=>x"8104",	-- 1000000100000100  brine	r0, fact_16.overflow
  589=>x"022E",	-- 0000001000101110  
  590=>x"0612",	-- 0000011000010010  dec	r2, r2
  591=>x"BE94",	-- 1011111010010100  brine	r2, fact_16.loop
  592=>x"E383",	-- 1110001110000011  ba	-, r6
  593=>x"063F",	-- 0000011000111111  dec	r7, r7
  594=>x"D23E",	-- 1101001000111110  sw	r6, r7
  595=>x"D013",	-- 1101000000010011  lw	r3, r2
  596=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  597=>x"84D8",	-- 1000010011011000  brieq	r3, puts.end
  598=>x"063F",	-- 0000011000111111  dec	r7, r7
  599=>x"D23A",	-- 1101001000111010  sw	r2, r7
  600=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  601=>x"026B",	-- 0000001001101011  
  602=>x"D03A",	-- 1101000000111010  lw	r2, r7
  603=>x"043F",	-- 0000010000111111  inc	r7, r7
  604=>x"D013",	-- 1101000000010011  lw	r3, r2
  605=>x"4E1B",	-- 0100111000011011  shl	r3, r3, 7
  606=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  607=>x"8258",	-- 1000001001011000  brieq	r3, puts.end
  608=>x"063F",	-- 0000011000111111  dec	r7, r7
  609=>x"D23A",	-- 1101001000111010  sw	r2, r7
  610=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  611=>x"026B",	-- 0000001001101011  
  612=>x"D03A",	-- 1101000000111010  lw	r2, r7
  613=>x"043F",	-- 0000010000111111  inc	r7, r7
  614=>x"0412",	-- 0000010000010010  inc	r2, r2
  615=>x"BB03",	-- 1011101100000011  bri	-, puts.loop
  616=>x"D03E",	-- 1101000000111110  lw	r6, r7
  617=>x"043F",	-- 0000010000111111  inc	r7, r7
  618=>x"E383",	-- 1110001110000011  ba	-, r6
  619=>x"063F",	-- 0000011000111111  dec	r7, r7
  620=>x"D23E",	-- 1101001000111110  sw	r6, r7
  621=>x"063F",	-- 0000011000111111  dec	r7, r7
  622=>x"D238",	-- 1101001000111000  sw	r0, r7
  623=>x"063F",	-- 0000011000111111  dec	r7, r7
  624=>x"D239",	-- 1101001000111001  sw	r1, r7
  625=>x"FFF2",	-- 1111111111110010  liw	r2, font_map
  626=>x"12C0",	-- 0001001011000000  
  627=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  628=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  629=>x"C043",	-- 1100000001000011  li	r3, 8
  630=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  631=>x"02D5",	-- 0000001011010101  
  632=>x"D039",	-- 1101000000111001  lw	r1, r7
  633=>x"043F",	-- 0000010000111111  inc	r7, r7
  634=>x"D038",	-- 1101000000111000  lw	r0, r7
  635=>x"043F",	-- 0000010000111111  inc	r7, r7
  636=>x"0400",	-- 0000010000000000  inc	r0, r0
  637=>x"D03E",	-- 1101000000111110  lw	r6, r7
  638=>x"043F",	-- 0000010000111111  inc	r7, r7
  639=>x"E383",	-- 1110001110000011  ba	-, r6
  640=>x"063F",	-- 0000011000111111  dec	r7, r7
  641=>x"D23E",	-- 1101001000111110  sw	r6, r7
  642=>x"FFF4",	-- 1111111111110100  liw	r4, 10000
  643=>x"2710",	-- 0010011100010000  
  644=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  645=>x"0293",	-- 0000001010010011  
  646=>x"FFF4",	-- 1111111111110100  liw	r4, 1000
  647=>x"03E8",	-- 0000001111101000  
  648=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  649=>x"0293",	-- 0000001010010011  
  650=>x"C324",	-- 1100001100100100  li	r4, 100
  651=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  652=>x"0293",	-- 0000001010010011  
  653=>x"C054",	-- 1100000001010100  li	r4, 10
  654=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  655=>x"0293",	-- 0000001010010011  
  656=>x"D03E",	-- 1101000000111110  lw	r6, r7
  657=>x"043F",	-- 0000010000111111  inc	r7, r7
  658=>x"C00C",	-- 1100000000001100  li	r4, 1
  659=>x"C17B",	-- 1100000101111011  li	r3, 0x2F
  660=>x"041B",	-- 0000010000011011  inc	r3, r3
  661=>x"0B12",	-- 0000101100010010  sub	r2, r2, r4
  662=>x"BF91",	-- 1011111110010001  brige	r2, printnum.loop
  663=>x"0912",	-- 0000100100010010  add	r2, r2, r4
  664=>x"063F",	-- 0000011000111111  dec	r7, r7
  665=>x"D23E",	-- 1101001000111110  sw	r6, r7
  666=>x"063F",	-- 0000011000111111  dec	r7, r7
  667=>x"D23A",	-- 1101001000111010  sw	r2, r7
  668=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  669=>x"026B",	-- 0000001001101011  
  670=>x"D03A",	-- 1101000000111010  lw	r2, r7
  671=>x"043F",	-- 0000010000111111  inc	r7, r7
  672=>x"D03E",	-- 1101000000111110  lw	r6, r7
  673=>x"043F",	-- 0000010000111111  inc	r7, r7
  674=>x"E383",	-- 1110001110000011  ba	-, r6
  675=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  676=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  677=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  678=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  679=>x"C0A0",	-- 1100000010100000  li	r0, 20
  680=>x"D011",	-- 1101000000010001  lw	r1, r2
  681=>x"D221",	-- 1101001000100001  sw	r1, r4
  682=>x"0412",	-- 0000010000010010  inc	r2, r2
  683=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  684=>x"061B",	-- 0000011000011011  dec	r3, r3
  685=>x"BEDC",	-- 1011111011011100  brine	r3, put_sprite_16_aligned.loop
  686=>x"E383",	-- 1110001110000011  ba	-, r6
  687=>x"C07D",	-- 1100000001111101  li	r5, 15
  688=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  689=>x"6600",	-- 0110011000000000  shr	r0, r0, 3
  690=>x"BC68",	-- 1011110001101000  brieq	r5, put_sprite_16_aligned
  691=>x"062D",	-- 0000011000101101  dec	r5, r5
  692=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  693=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  694=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  695=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  696=>x"063F",	-- 0000011000111111  dec	r7, r7
  697=>x"D23B",	-- 1101001000111011  sw	r3, r7
  698=>x"D011",	-- 1101000000010001  lw	r1, r2
  699=>x"CFF8",	-- 1100111111111000  li	r0, -1
  700=>x"3D40",	-- 0011110101000000  rsr	r0, r0, r5
  701=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  702=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  703=>x"D023",	-- 1101000000100011  lw	r3, r4
  704=>x"2600",	-- 0010011000000000  not	r0, r0
  705=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  706=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  707=>x"D221",	-- 1101001000100001  sw	r1, r4
  708=>x"0424",	-- 0000010000100100  inc	r4, r4
  709=>x"D011",	-- 1101000000010001  lw	r1, r2
  710=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  711=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  712=>x"D023",	-- 1101000000100011  lw	r3, r4
  713=>x"2600",	-- 0010011000000000  not	r0, r0
  714=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  715=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  716=>x"D221",	-- 1101001000100001  sw	r1, r4
  717=>x"0412",	-- 0000010000010010  inc	r2, r2
  718=>x"C098",	-- 1100000010011000  li	r0, 19
  719=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  720=>x"D03B",	-- 1101000000111011  lw	r3, r7
  721=>x"043F",	-- 0000010000111111  inc	r7, r7
  722=>x"061B",	-- 0000011000011011  dec	r3, r3
  723=>x"B95C",	-- 1011100101011100  brine	r3, put_sprite_16.loop
  724=>x"E383",	-- 1110001110000011  ba	-, r6
  725=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  726=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  727=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  728=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  729=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  730=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  731=>x"C0A5",	-- 1100000010100101  li	r5, 20
  732=>x"8404",	-- 1000010000000100  brine	r0, put_sprite_8_aligned.loop1
  733=>x"D010",	-- 1101000000010000  lw	r0, r2
  734=>x"D021",	-- 1101000000100001  lw	r1, r4
  735=>x"1A41",	-- 0001101001000001  mixhl	r1, r0, r1
  736=>x"D221",	-- 1101001000100001  sw	r1, r4
  737=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  738=>x"061B",	-- 0000011000011011  dec	r3, r3
  739=>x"E398",	-- 1110001110011000  baeq	r3, r6
  740=>x"D021",	-- 1101000000100001  lw	r1, r4
  741=>x"1E41",	-- 0001111001000001  mixll	r1, r0, r1
  742=>x"D221",	-- 1101001000100001  sw	r1, r4
  743=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  744=>x"0412",	-- 0000010000010010  inc	r2, r2
  745=>x"061B",	-- 0000011000011011  dec	r3, r3
  746=>x"E398",	-- 1110001110011000  baeq	r3, r6
  747=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop0
  748=>x"D010",	-- 1101000000010000  lw	r0, r2
  749=>x"D021",	-- 1101000000100001  lw	r1, r4
  750=>x"1809",	-- 0001100000001001  mixhh	r1, r1, r0
  751=>x"D221",	-- 1101001000100001  sw	r1, r4
  752=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  753=>x"061B",	-- 0000011000011011  dec	r3, r3
  754=>x"E398",	-- 1110001110011000  baeq	r3, r6
  755=>x"D021",	-- 1101000000100001  lw	r1, r4
  756=>x"1A09",	-- 0001101000001001  mixhl	r1, r1, r0
  757=>x"D221",	-- 1101001000100001  sw	r1, r4
  758=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  759=>x"0412",	-- 0000010000010010  inc	r2, r2
  760=>x"061B",	-- 0000011000011011  dec	r3, r3
  761=>x"E398",	-- 1110001110011000  baeq	r3, r6
  762=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop1
  763=>x"C03D",	-- 1100000000111101  li	r5, 7
  764=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  765=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  766=>x"B5E8",	-- 1011010111101000  brieq	r5, put_sprite_8_aligned
  767=>x"062D",	-- 0000011000101101  dec	r5, r5
  768=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  769=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  770=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  771=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  772=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  773=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  774=>x"8A04",	-- 1000101000000100  brine	r0, put_sprite_8.loop1
  775=>x"D010",	-- 1101000000010000  lw	r0, r2
  776=>x"063F",	-- 0000011000111111  dec	r7, r7
  777=>x"D23A",	-- 1101001000111010  sw	r2, r7
  778=>x"C802",	-- 1100100000000010  li	r2, 0x100
  779=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  780=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  781=>x"D021",	-- 1101000000100001  lw	r1, r4
  782=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  783=>x"2612",	-- 0010011000010010  not	r2, r2
  784=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  785=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  786=>x"D221",	-- 1101001000100001  sw	r1, r4
  787=>x"C0A1",	-- 1100000010100001  li	r1, 20
  788=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  789=>x"D03A",	-- 1101000000111010  lw	r2, r7
  790=>x"043F",	-- 0000010000111111  inc	r7, r7
  791=>x"061B",	-- 0000011000011011  dec	r3, r3
  792=>x"E398",	-- 1110001110011000  baeq	r3, r6
  793=>x"D010",	-- 1101000000010000  lw	r0, r2
  794=>x"063F",	-- 0000011000111111  dec	r7, r7
  795=>x"D23A",	-- 1101001000111010  sw	r2, r7
  796=>x"1E00",	-- 0001111000000000  mixll	r0, r0, r0
  797=>x"C802",	-- 1100100000000010  li	r2, 0x100
  798=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  799=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  800=>x"D021",	-- 1101000000100001  lw	r1, r4
  801=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  802=>x"2612",	-- 0010011000010010  not	r2, r2
  803=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  804=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  805=>x"D221",	-- 1101001000100001  sw	r1, r4
  806=>x"C0A1",	-- 1100000010100001  li	r1, 20
  807=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  808=>x"D03A",	-- 1101000000111010  lw	r2, r7
  809=>x"043F",	-- 0000010000111111  inc	r7, r7
  810=>x"0412",	-- 0000010000010010  inc	r2, r2
  811=>x"061B",	-- 0000011000011011  dec	r3, r3
  812=>x"E398",	-- 1110001110011000  baeq	r3, r6
  813=>x"B683",	-- 1011011010000011  bri	-, put_sprite_8.loop0
  814=>x"D010",	-- 1101000000010000  lw	r0, r2
  815=>x"063F",	-- 0000011000111111  dec	r7, r7
  816=>x"D23A",	-- 1101001000111010  sw	r2, r7
  817=>x"063F",	-- 0000011000111111  dec	r7, r7
  818=>x"D23B",	-- 1101001000111011  sw	r3, r7
  819=>x"C802",	-- 1100100000000010  li	r2, 0x100
  820=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  821=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  822=>x"2080",	-- 0010000010000000  and	r0, r0, r2
  823=>x"D021",	-- 1101000000100001  lw	r1, r4
  824=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
  825=>x"261B",	-- 0010011000011011  not	r3, r3
  826=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  827=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
  828=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  829=>x"D221",	-- 1101001000100001  sw	r1, r4
  830=>x"0424",	-- 0000010000100100  inc	r4, r4
  831=>x"D021",	-- 1101000000100001  lw	r1, r4
  832=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  833=>x"261B",	-- 0010011000011011  not	r3, r3
  834=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  835=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
  836=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  837=>x"D221",	-- 1101001000100001  sw	r1, r4
  838=>x"C099",	-- 1100000010011001  li	r1, 19
  839=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  840=>x"D03B",	-- 1101000000111011  lw	r3, r7
  841=>x"043F",	-- 0000010000111111  inc	r7, r7
  842=>x"D03A",	-- 1101000000111010  lw	r2, r7
  843=>x"043F",	-- 0000010000111111  inc	r7, r7
  844=>x"061B",	-- 0000011000011011  dec	r3, r3
  845=>x"E398",	-- 1110001110011000  baeq	r3, r6
  846=>x"D010",	-- 1101000000010000  lw	r0, r2
  847=>x"4E00",	-- 0100111000000000  shl	r0, r0, 7
  848=>x"063F",	-- 0000011000111111  dec	r7, r7
  849=>x"D23A",	-- 1101001000111010  sw	r2, r7
  850=>x"063F",	-- 0000011000111111  dec	r7, r7
  851=>x"D23B",	-- 1101001000111011  sw	r3, r7
  852=>x"C802",	-- 1100100000000010  li	r2, 0x100
  853=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  854=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  855=>x"2080",	-- 0010000010000000  and	r0, r0, r2
  856=>x"D021",	-- 1101000000100001  lw	r1, r4
  857=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
  858=>x"261B",	-- 0010011000011011  not	r3, r3
  859=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  860=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
  861=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  862=>x"D221",	-- 1101001000100001  sw	r1, r4
  863=>x"0424",	-- 0000010000100100  inc	r4, r4
  864=>x"D021",	-- 1101000000100001  lw	r1, r4
  865=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  866=>x"261B",	-- 0010011000011011  not	r3, r3
  867=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  868=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
  869=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  870=>x"D221",	-- 1101001000100001  sw	r1, r4
  871=>x"C099",	-- 1100000010011001  li	r1, 19
  872=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  873=>x"D03B",	-- 1101000000111011  lw	r3, r7
  874=>x"043F",	-- 0000010000111111  inc	r7, r7
  875=>x"D03A",	-- 1101000000111010  lw	r2, r7
  876=>x"043F",	-- 0000010000111111  inc	r7, r7
  877=>x"0412",	-- 0000010000010010  inc	r2, r2
  878=>x"061B",	-- 0000011000011011  dec	r3, r3
  879=>x"E398",	-- 1110001110011000  baeq	r3, r6
  880=>x"AF83",	-- 1010111110000011  bri	-, put_sprite_8.loop1
    others => x"0000"
    );
begin
  process(CLK)
  begin
    if (CLK'event AND CLK='1') then
      D <= m(to_integer(unsigned(AD)));
    end if;
  end process;
end Behavioral;
