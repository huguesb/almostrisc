----------------------------------------------------------------------------------
--
-- File retrieved, on 07/02/2010, from :
-- http://sebastien-viardot.imag.fr/Enseignements/Archi1A2s/sources/ROMPROG.vhd
--
-- Slightly altered to get rid of vendor-specific packages and adjust formatting
-- Now auto-filled by asrom script
--
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROMPROG is
  Port ( AD : in  STD_LOGIC_VECTOR (12 downto 0);
         D : out  STD_LOGIC_VECTOR (15 downto 0);
         CLK : in STD_LOGIC);
end ROMPROG;

architecture Behavioral of ROMPROG is
  constant low_address: natural := 0;
  constant high_address: natural := 8192;
  subtype octet is std_logic_vector( 15 downto 0 );
  type zone_memoire is
    array (natural range low_address to high_address-1) of octet;
  constant m: zone_memoire:= (
    0=>x"FFF7",	-- 1111111111110111  liw	r7, IRQ_mask
    1=>x"2000",	-- 0010000000000000  
    2=>x"F8C0",	-- 1111100011000000  bai	-, os_init
    3=>x"0100",	-- 0000000100000000  
   16=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_ack
   17=>x"2002",	-- 0010000000000010  
   18=>x"D001",	-- 1101000000000001  lw	r1, r0
   19=>x"F54A",	-- 1111010101001010  bspl	r2, r1, 5
   20=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_error
   21=>x"0050",	-- 0000000001010000  
   22=>x"F4CA",	-- 1111010011001010  bspl	r2, r1, 3
   23=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_kbd
   24=>x"0060",	-- 0000000001100000  
   25=>x"F40A",	-- 1111010000001010  bspl	r2, r1, 0
   26=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_tmr
   27=>x"0040",	-- 0000000001000000  
   28=>x"D201",	-- 1101001000000001  sw	r1, r0
   29=>x"FFFE",	-- 1111111111111110  reti
   64=>x"263F",	-- 0010011000111111  not r7, r7
   65=>x"D7C0",	-- 1101011111000000  out	r7
   66=>x"E383",	-- 1110001110000011  ba	-, r6
   80=>x"25FF",	-- 0010010111111111  xor	r7, r7, r7
   81=>x"D7C0",	-- 1101011111000000  out	r7
   82=>x"E383",	-- 1110001110000011  ba	-, r6
   96=>x"FFF2",	-- 1111111111110010  liw	r2, PS2_rx
   97=>x"2004",	-- 0010000000000100  
   98=>x"D012",	-- 1101000000010010  lw	r2, r2
   99=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map + 8
  100=>x"1808",	-- 0001100000001000  
  101=>x"D01B",	-- 1101000000011011  lw	r3, r3
  102=>x"1EBF",	-- 0001111010111111  mixll	r7, r7, r2
  103=>x"C784",	-- 1100011110000100  li	r4, 0xF0
  104=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  105=>x"8B20",	-- 1000101100100000  brieq	r4, int_kbd.release
  106=>x"C704",	-- 1100011100000100  li	r4, 0xE0
  107=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  108=>x"88E0",	-- 1000100011100000  brieq	r4, int_kbd.extended
  109=>x"FFF5",	-- 1111111111110101  liw	r5, 0x16C0 - 1
  110=>x"16BF",	-- 0001011010111111  
  111=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  112=>x"80E0",	-- 1000000011100000  brieq	r4, $+3
  113=>x"FFF5",	-- 1111111111110101  liw	r5, 0x16CA - 1
  114=>x"16C9",	-- 0001011011001001  
  115=>x"042D",	-- 0000010000101101  inc	r5, r5
  116=>x"D02C",	-- 1101000000101100  lw	r4, r5
  117=>x"8560",	-- 1000010101100000  brieq	r4, scan_code_mismatch
  118=>x"6E24",	-- 0110111000100100  shr	r4, r4, 7
  119=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  120=>x"BEE4",	-- 1011111011100100  brine	r4, scan_code_loop
  121=>x"D02A",	-- 1101000000101010  lw	r2, r5
  122=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  123=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  124=>x"741B",	-- 0111010000011011  shr	r3, r3, 10
  125=>x"C00D",	-- 1100000000001101  li	r5, 1
  126=>x"0612",	-- 0000011000010010  dec	r2, r2
  127=>x"3AAA",	-- 0011101010101010  rrl	r2, r5, r2
  128=>x"FFF5",	-- 1111111111110101  liw	r5, key_press_map
  129=>x"1800",	-- 0001100000000000  
  130=>x"08ED",	-- 0000100011101101  add	r5, r5, r3
  131=>x"D02B",	-- 1101000000101011  lw	r3, r5
  132=>x"80E4",	-- 1000000011100100  brine	r4, scan_code_release
  133=>x"229B",	-- 0010001010011011  or	r3, r3, r2
  134=>x"80C3",	-- 1000000011000011  bri	-, scan_code_notify
  135=>x"2612",	-- 0010011000010010  not	r2, r2
  136=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  137=>x"D22B",	-- 1101001000101011  sw	r3, r5
  138=>x"C003",	-- 1100000000000011  li	r3, 0
  139=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  140=>x"1808",	-- 0001100000001000  
  141=>x"D223",	-- 1101001000100011  sw	r3, r4
  142=>x"E383",	-- 1110001110000011  ba	-, r6
  143=>x"C014",	-- 1100000000010100  li	r4, 2
  144=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  145=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  146=>x"1808",	-- 0001100000001000  
  147=>x"D223",	-- 1101001000100011  sw	r3, r4
  148=>x"E383",	-- 1110001110000011  ba	-, r6
  149=>x"C00C",	-- 1100000000001100  li	r4, 1
  150=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  151=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  152=>x"1808",	-- 0001100000001000  
  153=>x"D223",	-- 1101001000100011  sw	r3, r4
  154=>x"E383",	-- 1110001110000011  ba	-, r6
  256=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_mask
  257=>x"2000",	-- 0010000000000000  
  258=>x"C0C9",	-- 1100000011001001  li	r1, 0x19
  259=>x"D201",	-- 1101001000000001  sw	r1, r0
  260=>x"0400",	-- 0000010000000000  inc	r0, r0
  261=>x"CFF9",	-- 1100111111111001  li	r1, -1
  262=>x"D201",	-- 1101001000000001  sw	r1, r0
  263=>x"C03A",	-- 1100000000111010  li	r2, 7
  264=>x"0880",	-- 0000100010000000  add	r0, r0, r2
  265=>x"C0EA",	-- 1100000011101010  li	r2, 0x1D
  266=>x"D202",	-- 1101001000000010  sw	r2, r0
  267=>x"0400",	-- 0000010000000000  inc	r0, r0
  268=>x"C07A",	-- 1100000001111010  li	r2, 15
  269=>x"D202",	-- 1101001000000010  sw	r2, r0
  270=>x"FFF0",	-- 1111111111110000  liw	r0, key_press_map
  271=>x"1800",	-- 0001100000000000  
  272=>x"C001",	-- 1100000000000001  li	r1, 0
  273=>x"C042",	-- 1100000001000010  li	r2, 8
  274=>x"D201",	-- 1101001000000001  sw	r1, r0
  275=>x"0400",	-- 0000010000000000  inc	r0, r0
  276=>x"0612",	-- 0000011000010010  dec	r2, r2
  277=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  278=>x"C0F3",	-- 1100000011110011  li	r3, 30
  279=>x"CFFA",	-- 1100111111111010  li	r2, -1
  280=>x"D21A",	-- 1101001000011010  sw	r2, r3
  281=>x"8083",	-- 1000000010000011  bri	-, PaperGameStart
  282=>x"8003",	-- 1000000000000011  bri	-, PaperMenuLoop
  283=>x"C000",	-- 1100000000000000  li	r0, 0
  284=>x"FFF1",	-- 1111111111110001  liw	r1, 0x0801
  285=>x"0801",	-- 0000100000000001  
  286=>x"063F",	-- 0000011000111111  dec	r7, r7
  287=>x"D238",	-- 1101001000111000  sw	r0, r7
  288=>x"063F",	-- 0000011000111111  dec	r7, r7
  289=>x"D239",	-- 1101001000111001  sw	r1, r7
  290=>x"063F",	-- 0000011000111111  dec	r7, r7
  291=>x"D23A",	-- 1101001000111010  sw	r2, r7
  292=>x"C000",	-- 1100000000000000  li	r0, 0
  293=>x"CFF9",	-- 1100111111111001  li	r1, -1
  294=>x"C0A2",	-- 1100000010100010  li	r2, 20
  295=>x"D201",	-- 1101001000000001  sw	r1, r0
  296=>x"0400",	-- 0000010000000000  inc	r0, r0
  297=>x"0612",	-- 0000011000010010  dec	r2, r2
  298=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  299=>x"C001",	-- 1100000000000001  li	r1, 0
  300=>x"FFF2",	-- 1111111111110010  liw	r2, 18*20
  301=>x"0168",	-- 0000000101101000  
  302=>x"D201",	-- 1101001000000001  sw	r1, r0
  303=>x"0400",	-- 0000010000000000  inc	r0, r0
  304=>x"0612",	-- 0000011000010010  dec	r2, r2
  305=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  306=>x"CFF9",	-- 1100111111111001  li	r1, -1
  307=>x"C0A2",	-- 1100000010100010  li	r2, 20
  308=>x"D201",	-- 1101001000000001  sw	r1, r0
  309=>x"0400",	-- 0000010000000000  inc	r0, r0
  310=>x"0612",	-- 0000011000010010  dec	r2, r2
  311=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  312=>x"C020",	-- 1100000000100000  li	r0, 4
  313=>x"C029",	-- 1100000000101001  li	r1, 5
  314=>x"FFF2",	-- 1111111111110010  liw	r2, paper_title
  315=>x"1730",	-- 0001011100110000  
  316=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  317=>x"0200",	-- 0000001000000000  
  318=>x"C790",	-- 1100011110010000  li	r0, 242
  319=>x"C009",	-- 1100000000001001  li	r1, 1
  320=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud
  321=>x"1720",	-- 0001011100100000  
  322=>x"C043",	-- 1100000001000011  li	r3, 8
  323=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  324=>x"028B",	-- 0000001010001011  
  325=>x"C118",	-- 1100000100011000  li	r0, 35
  326=>x"C009",	-- 1100000000001001  li	r1, 1
  327=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  328=>x"1736",	-- 0001011100110110  
  329=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  330=>x"0200",	-- 0000001000000000  
  331=>x"C790",	-- 1100011110010000  li	r0, 242
  332=>x"C051",	-- 1100000001010001  li	r1, 10
  333=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud + 4
  334=>x"1724",	-- 0001011100100100  
  335=>x"C043",	-- 1100000001000011  li	r3, 8
  336=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  337=>x"028B",	-- 0000001010001011  
  338=>x"C118",	-- 1100000100011000  li	r0, 35
  339=>x"C051",	-- 1100000001010001  li	r1, 10
  340=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  341=>x"1736",	-- 0001011100110110  
  342=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  343=>x"0200",	-- 0000001000000000  
  344=>x"D03A",	-- 1101000000111010  lw	r2, r7
  345=>x"043F",	-- 0000010000111111  inc	r7, r7
  346=>x"D039",	-- 1101000000111001  lw	r1, r7
  347=>x"043F",	-- 0000010000111111  inc	r7, r7
  348=>x"D038",	-- 1101000000111000  lw	r0, r7
  349=>x"043F",	-- 0000010000111111  inc	r7, r7
  350=>x"063F",	-- 0000011000111111  dec	r7, r7
  351=>x"D238",	-- 1101001000111000  sw	r0, r7
  352=>x"063F",	-- 0000011000111111  dec	r7, r7
  353=>x"D239",	-- 1101001000111001  sw	r1, r7
  354=>x"063F",	-- 0000011000111111  dec	r7, r7
  355=>x"D23A",	-- 1101001000111010  sw	r2, r7
  356=>x"CC80",	-- 1100110010000000  li	r0, 20*20
  357=>x"C001",	-- 1100000000000001  li	r1, 0
  358=>x"FFF2",	-- 1111111111110010  liw	r2, 220*20
  359=>x"1130",	-- 0001000100110000  
  360=>x"D201",	-- 1101001000000001  sw	r1, r0
  361=>x"0400",	-- 0000010000000000  inc	r0, r0
  362=>x"0612",	-- 0000011000010010  dec	r2, r2
  363=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  364=>x"C4C0",	-- 1100010011000000  li	r0, 152
  365=>x"C161",	-- 1100000101100001  li	r1, 44
  366=>x"FFF2",	-- 1111111111110010  liw	r2, paper_sprites
  367=>x"16D0",	-- 0001011011010000  
  368=>x"C083",	-- 1100000010000011  li	r3, 16
  369=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_16
  370=>x"023B",	-- 0000001000111011  
  371=>x"D03A",	-- 1101000000111010  lw	r2, r7
  372=>x"043F",	-- 0000010000111111  inc	r7, r7
  373=>x"D039",	-- 1101000000111001  lw	r1, r7
  374=>x"043F",	-- 0000010000111111  inc	r7, r7
  375=>x"D038",	-- 1101000000111000  lw	r0, r7
  376=>x"043F",	-- 0000010000111111  inc	r7, r7
  377=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  378=>x"1800",	-- 0001100000000000  
  379=>x"D01B",	-- 1101000000011011  lw	r3, r3
  380=>x"9518",	-- 1001010100011000  brieq	r3, event_not_kbd
  381=>x"F7DC",	-- 1111011111011100  bspl	r4, r3, 15
  382=>x"82A0",	-- 1000001010100000  brieq	r4, PaperGameQuit
  383=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  384=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveUp
  385=>x"F49C",	-- 1111010010011100  bspl	r4, r3, 2
  386=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveDOWN
  387=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  388=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveLEFT
  389=>x"F4DC",	-- 1111010011011100  bspl	r4, r3, 3
  390=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveRIGHT
  391=>x"BC83",	-- 1011110010000011  bri	-, PaperGameLoop
  392=>x"FFFF",	-- 1111111111111111  reset
  393=>x"C040",	-- 1100000001000000  li	r0, 8
  394=>x"C041",	-- 1100000001000001  li	r1, 8
  395=>x"063F",	-- 0000011000111111  dec	r7, r7
  396=>x"D239",	-- 1101001000111001  sw	r1, r7
  397=>x"063F",	-- 0000011000111111  dec	r7, r7
  398=>x"D238",	-- 1101001000111000  sw	r0, r7
  399=>x"FFF2",	-- 1111111111110010  liw	r2, font_map + 4 * 0x23
  400=>x"134C",	-- 0001001101001100  
  401=>x"C043",	-- 1100000001000011  li	r3, 8
  402=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  403=>x"028B",	-- 0000001010001011  
  404=>x"D038",	-- 1101000000111000  lw	r0, r7
  405=>x"043F",	-- 0000010000111111  inc	r7, r7
  406=>x"D039",	-- 1101000000111001  lw	r1, r7
  407=>x"043F",	-- 0000010000111111  inc	r7, r7
  408=>x"C0A2",	-- 1100000010100010  li	r2, 20
  409=>x"C003",	-- 1100000000000011  li	r3, 0
  410=>x"061B",	-- 0000011000011011  dec	r3, r3
  411=>x"BFDC",	-- 1011111111011100  brine	r3, $-1
  412=>x"0612",	-- 0000011000010010  dec	r2, r2
  413=>x"BF14",	-- 1011111100010100  brine	r2, $-4
  414=>x"FFF2",	-- 1111111111110010  liw	r2, key_press_map
  415=>x"1800",	-- 0001100000000000  
  416=>x"D012",	-- 1101000000010010  lw	r2, r2
  417=>x"8BD0",	-- 1000101111010000  brieq	r2, event_not_kbd
  418=>x"063F",	-- 0000011000111111  dec	r7, r7
  419=>x"D23A",	-- 1101001000111010  sw	r2, r7
  420=>x"063F",	-- 0000011000111111  dec	r7, r7
  421=>x"D239",	-- 1101001000111001  sw	r1, r7
  422=>x"063F",	-- 0000011000111111  dec	r7, r7
  423=>x"D238",	-- 1101001000111000  sw	r0, r7
  424=>x"FFF2",	-- 1111111111110010  liw	r2, font_map
  425=>x"12C0",	-- 0001001011000000  
  426=>x"C043",	-- 1100000001000011  li	r3, 8
  427=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  428=>x"028B",	-- 0000001010001011  
  429=>x"D038",	-- 1101000000111000  lw	r0, r7
  430=>x"043F",	-- 0000010000111111  inc	r7, r7
  431=>x"D039",	-- 1101000000111001  lw	r1, r7
  432=>x"043F",	-- 0000010000111111  inc	r7, r7
  433=>x"D03A",	-- 1101000000111010  lw	r2, r7
  434=>x"043F",	-- 0000010000111111  inc	r7, r7
  435=>x"F413",	-- 1111010000010011  bspl	r3, r2, 0
  436=>x"81D8",	-- 1000000111011000  brieq	r3, event_kbd_no_up
  437=>x"C043",	-- 1100000001000011  li	r3, 8
  438=>x"0ACB",	-- 0000101011001011  sub	r3, r1, r3
  439=>x"809C",	-- 1000000010011100  brine	r3, event_kbd_no_clip_up
  440=>x"C781",	-- 1100011110000001  li	r1, 240
  441=>x"C043",	-- 1100000001000011  li	r3, 8
  442=>x"0AC9",	-- 0000101011001001  sub	r1, r1, r3
  443=>x"F453",	-- 1111010001010011  bspl	r3, r2, 1
  444=>x"8118",	-- 1000000100011000  brieq	r3, event_kbd_no_left
  445=>x"8084",	-- 1000000010000100  brine	r0, event_kbd_no_clip_left
  446=>x"C9C0",	-- 1100100111000000  li	r0, 39*8
  447=>x"0600",	-- 0000011000000000  dec	r0, r0
  448=>x"F493",	-- 1111010010010011  bspl	r3, r2, 2
  449=>x"81D8",	-- 1000000111011000  brieq	r3, event_kbd_no_down
  450=>x"C743",	-- 1100011101000011  li	r3, 232
  451=>x"0ACB",	-- 0000101011001011  sub	r3, r1, r3
  452=>x"809D",	-- 1000000010011101  brilt	r3, event_kbd_no_clip_down
  453=>x"C001",	-- 1100000000000001  li	r1, 0
  454=>x"C043",	-- 1100000001000011  li	r3, 8
  455=>x"08C9",	-- 0000100011001001  add	r1, r1, r3
  456=>x"F4D3",	-- 1111010011010011  bspl	r3, r2, 3
  457=>x"8198",	-- 1000000110011000  brieq	r3, event_kbd_no_right
  458=>x"C9C3",	-- 1100100111000011  li	r3, 39*8
  459=>x"0AC3",	-- 0000101011000011  sub	r3, r0, r3
  460=>x"809D",	-- 1000000010011101  brilt	r3, event_kbd_no_clip_right
  461=>x"CFF8",	-- 1100111111111000  li	r0, -1
  462=>x"0400",	-- 0000010000000000  inc	r0, r0
  463=>x"AF03",	-- 1010111100000011  bri	-, redraw
  464=>x"B383",	-- 1011001110000011  bri	-, event_loop
  465=>x"C750",	-- 1100011101010000  li	r0, 234
  466=>x"C1C2",	-- 1100000111000010  li	r2, 56
  467=>x"FAC6",	-- 1111101011000110  bail	-, r6, div_16_16
  468=>x"01E9",	-- 0000000111101001  
  469=>x"C448",	-- 1100010001001000  li	r0, 137
  470=>x"C472",	-- 1100010001110010  li	r2, 142
  471=>x"FAC6",	-- 1111101011000110  bail	-, r6, mult_16_16
  472=>x"01DD",	-- 0000000111011101  
  473=>x"C03A",	-- 1100000000111010  li r2, 7
  474=>x"FAC6",	-- 1111101011000110  bail	-, r6, fact_16
  475=>x"01F4",	-- 0000000111110100  
  476=>x"FFFF",	-- 1111111111111111  reset
  477=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  478=>x"2524",	-- 0010010100100100  xor	r4, r4, r4
  479=>x"C085",	-- 1100000010000101  li	r5, 16
  480=>x"0849",	-- 0000100001001001  add	r1, r1, r1
  481=>x"0C00",	-- 0000110000000000  adc	r0, r0, r0
  482=>x"0EDB",	-- 0000111011011011  sbc	r3, r3, r3
  483=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  484=>x"08C9",	-- 0000100011001001  add	r1, r1, r3
  485=>x"0D00",	-- 0000110100000000  adc	r0, r0, r4
  486=>x"062D",	-- 0000011000101101  dec	r5, r5
  487=>x"BE6C",	-- 1011111001101100  brine	r5, mult_16_16.loop
  488=>x"E383",	-- 1110001110000011  ba	-, r6
  489=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  490=>x"C084",	-- 1100000010000100  li	r4, 16
  491=>x"0800",	-- 0000100000000000  add	r0, r0, r0
  492=>x"0C49",	-- 0000110001001001  adc	r1, r1, r1
  493=>x"0A8B",	-- 0000101010001011  sub	r3, r1, r2
  494=>x"80DD",	-- 1000000011011101  brilt	r3, div_16_16.skip
  495=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  496=>x"0400",	-- 0000010000000000  inc	r0, r0
  497=>x"0624",	-- 0000011000100100  dec	r4, r4
  498=>x"BE64",	-- 1011111001100100  brine	r4, div_16_16.loop
  499=>x"E383",	-- 1110001110000011  ba	-, r6
  500=>x"2400",	-- 0010010000000000  xor	r0, r0, r0
  501=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  502=>x"8250",	-- 1000001001010000  brieq	r2, fact_16.end
  503=>x"0409",	-- 0000010000001001  inc	r1, r1
  504=>x"1008",	-- 0001000000001000  mova	r0, r1
  505=>x"FAC6",	-- 1111101011000110  bail	-, r6, mult_16_16
  506=>x"01DD",	-- 0000000111011101  
  507=>x"8104",	-- 1000000100000100  brine	r0, fact_16.overflow
  508=>x"01DD",	-- 0000000111011101  
  509=>x"0612",	-- 0000011000010010  dec	r2, r2
  510=>x"BE94",	-- 1011111010010100  brine	r2, fact_16.loop
  511=>x"E383",	-- 1110001110000011  ba	-, r6
  512=>x"063F",	-- 0000011000111111  dec	r7, r7
  513=>x"D23E",	-- 1101001000111110  sw	r6, r7
  514=>x"D013",	-- 1101000000010011  lw	r3, r2
  515=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  516=>x"84D8",	-- 1000010011011000  brieq	r3, puts.end
  517=>x"063F",	-- 0000011000111111  dec	r7, r7
  518=>x"D23A",	-- 1101001000111010  sw	r2, r7
  519=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  520=>x"021A",	-- 0000001000011010  
  521=>x"D03A",	-- 1101000000111010  lw	r2, r7
  522=>x"043F",	-- 0000010000111111  inc	r7, r7
  523=>x"D013",	-- 1101000000010011  lw	r3, r2
  524=>x"4E1B",	-- 0100111000011011  shl	r3, r3, 7
  525=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  526=>x"8258",	-- 1000001001011000  brieq	r3, puts.end
  527=>x"063F",	-- 0000011000111111  dec	r7, r7
  528=>x"D23A",	-- 1101001000111010  sw	r2, r7
  529=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  530=>x"021A",	-- 0000001000011010  
  531=>x"D03A",	-- 1101000000111010  lw	r2, r7
  532=>x"043F",	-- 0000010000111111  inc	r7, r7
  533=>x"0412",	-- 0000010000010010  inc	r2, r2
  534=>x"BB03",	-- 1011101100000011  bri	-, puts.loop
  535=>x"D03E",	-- 1101000000111110  lw	r6, r7
  536=>x"043F",	-- 0000010000111111  inc	r7, r7
  537=>x"E383",	-- 1110001110000011  ba	-, r6
  538=>x"063F",	-- 0000011000111111  dec	r7, r7
  539=>x"D23E",	-- 1101001000111110  sw	r6, r7
  540=>x"063F",	-- 0000011000111111  dec	r7, r7
  541=>x"D238",	-- 1101001000111000  sw	r0, r7
  542=>x"063F",	-- 0000011000111111  dec	r7, r7
  543=>x"D239",	-- 1101001000111001  sw	r1, r7
  544=>x"FFF2",	-- 1111111111110010  liw	r2, font_map
  545=>x"12C0",	-- 0001001011000000  
  546=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  547=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  548=>x"C043",	-- 1100000001000011  li	r3, 8
  549=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  550=>x"0265",	-- 0000001001100101  
  551=>x"D039",	-- 1101000000111001  lw	r1, r7
  552=>x"043F",	-- 0000010000111111  inc	r7, r7
  553=>x"D038",	-- 1101000000111000  lw	r0, r7
  554=>x"043F",	-- 0000010000111111  inc	r7, r7
  555=>x"0400",	-- 0000010000000000  inc	r0, r0
  556=>x"D03E",	-- 1101000000111110  lw	r6, r7
  557=>x"043F",	-- 0000010000111111  inc	r7, r7
  558=>x"E383",	-- 1110001110000011  ba	-, r6
  559=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  560=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  561=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  562=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  563=>x"C0A0",	-- 1100000010100000  li	r0, 20
  564=>x"D011",	-- 1101000000010001  lw	r1, r2
  565=>x"D221",	-- 1101001000100001  sw	r1, r4
  566=>x"0412",	-- 0000010000010010  inc	r2, r2
  567=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  568=>x"061B",	-- 0000011000011011  dec	r3, r3
  569=>x"BEDC",	-- 1011111011011100  brine	r3, put_sprite_16_aligned.loop
  570=>x"E383",	-- 1110001110000011  ba	-, r6
  571=>x"C07D",	-- 1100000001111101  li	r5, 15
  572=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  573=>x"6600",	-- 0110011000000000  shr	r0, r0, 3
  574=>x"BC68",	-- 1011110001101000  brieq	r5, put_sprite_16_aligned
  575=>x"062D",	-- 0000011000101101  dec	r5, r5
  576=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  577=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  578=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  579=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  580=>x"063F",	-- 0000011000111111  dec	r7, r7
  581=>x"D23B",	-- 1101001000111011  sw	r3, r7
  582=>x"D011",	-- 1101000000010001  lw	r1, r2
  583=>x"CFF8",	-- 1100111111111000  li	r0, -1
  584=>x"3D40",	-- 0011110101000000  rsr	r0, r0, r5
  585=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  586=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  587=>x"D023",	-- 1101000000100011  lw	r3, r4
  588=>x"2600",	-- 0010011000000000  not	r0, r0
  589=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  590=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  591=>x"D221",	-- 1101001000100001  sw	r1, r4
  592=>x"0424",	-- 0000010000100100  inc	r4, r4
  593=>x"D011",	-- 1101000000010001  lw	r1, r2
  594=>x"262D",	-- 0010011000101101  not	r5, r5
  595=>x"CFF8",	-- 1100111111111000  li	r0, -1
  596=>x"3F40",	-- 0011111101000000  rsl	r0, r0, r5
  597=>x"3B49",	-- 0011101101001001  rrl	r1, r1, r5
  598=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  599=>x"262D",	-- 0010011000101101  not	r5, r5
  600=>x"D023",	-- 1101000000100011  lw	r3, r4
  601=>x"2600",	-- 0010011000000000  not	r0, r0
  602=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  603=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  604=>x"D221",	-- 1101001000100001  sw	r1, r4
  605=>x"0412",	-- 0000010000010010  inc	r2, r2
  606=>x"C098",	-- 1100000010011000  li	r0, 19
  607=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  608=>x"D03B",	-- 1101000000111011  lw	r3, r7
  609=>x"043F",	-- 0000010000111111  inc	r7, r7
  610=>x"061B",	-- 0000011000011011  dec	r3, r3
  611=>x"B85C",	-- 1011100001011100  brine	r3, put_sprite_16.loop
  612=>x"E383",	-- 1110001110000011  ba	-, r6
  613=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  614=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  615=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  616=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  617=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  618=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  619=>x"C0A5",	-- 1100000010100101  li	r5, 20
  620=>x"8404",	-- 1000010000000100  brine	r0, put_sprite_8_aligned.loop1
  621=>x"D010",	-- 1101000000010000  lw	r0, r2
  622=>x"D021",	-- 1101000000100001  lw	r1, r4
  623=>x"1A41",	-- 0001101001000001  mixhl	r1, r0, r1
  624=>x"D221",	-- 1101001000100001  sw	r1, r4
  625=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  626=>x"061B",	-- 0000011000011011  dec	r3, r3
  627=>x"E398",	-- 1110001110011000  baeq	r3, r6
  628=>x"D021",	-- 1101000000100001  lw	r1, r4
  629=>x"1E41",	-- 0001111001000001  mixll	r1, r0, r1
  630=>x"D221",	-- 1101001000100001  sw	r1, r4
  631=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  632=>x"0412",	-- 0000010000010010  inc	r2, r2
  633=>x"061B",	-- 0000011000011011  dec	r3, r3
  634=>x"E398",	-- 1110001110011000  baeq	r3, r6
  635=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop0
  636=>x"D010",	-- 1101000000010000  lw	r0, r2
  637=>x"D021",	-- 1101000000100001  lw	r1, r4
  638=>x"1809",	-- 0001100000001001  mixhh	r1, r1, r0
  639=>x"D221",	-- 1101001000100001  sw	r1, r4
  640=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  641=>x"061B",	-- 0000011000011011  dec	r3, r3
  642=>x"E398",	-- 1110001110011000  baeq	r3, r6
  643=>x"D021",	-- 1101000000100001  lw	r1, r4
  644=>x"1A09",	-- 0001101000001001  mixhl	r1, r1, r0
  645=>x"D221",	-- 1101001000100001  sw	r1, r4
  646=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  647=>x"0412",	-- 0000010000010010  inc	r2, r2
  648=>x"061B",	-- 0000011000011011  dec	r3, r3
  649=>x"E398",	-- 1110001110011000  baeq	r3, r6
  650=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop1
  651=>x"C03D",	-- 1100000000111101  li	r5, 7
  652=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  653=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  654=>x"B5E8",	-- 1011010111101000  brieq	r5, put_sprite_8_aligned
  655=>x"062D",	-- 0000011000101101  dec	r5, r5
  656=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  657=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  658=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  659=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  660=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  661=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  662=>x"8A04",	-- 1000101000000100  brine	r0, put_sprite_8.loop1
  663=>x"D010",	-- 1101000000010000  lw	r0, r2
  664=>x"063F",	-- 0000011000111111  dec	r7, r7
  665=>x"D23A",	-- 1101001000111010  sw	r2, r7
  666=>x"C802",	-- 1100100000000010  li	r2, 0x100
  667=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  668=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  669=>x"D021",	-- 1101000000100001  lw	r1, r4
  670=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  671=>x"2612",	-- 0010011000010010  not	r2, r2
  672=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  673=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  674=>x"D221",	-- 1101001000100001  sw	r1, r4
  675=>x"C0A1",	-- 1100000010100001  li	r1, 20
  676=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  677=>x"D03A",	-- 1101000000111010  lw	r2, r7
  678=>x"043F",	-- 0000010000111111  inc	r7, r7
  679=>x"061B",	-- 0000011000011011  dec	r3, r3
  680=>x"E398",	-- 1110001110011000  baeq	r3, r6
  681=>x"D010",	-- 1101000000010000  lw	r0, r2
  682=>x"063F",	-- 0000011000111111  dec	r7, r7
  683=>x"D23A",	-- 1101001000111010  sw	r2, r7
  684=>x"1E00",	-- 0001111000000000  mixll	r0, r0, r0
  685=>x"C802",	-- 1100100000000010  li	r2, 0x100
  686=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  687=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  688=>x"D021",	-- 1101000000100001  lw	r1, r4
  689=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  690=>x"2612",	-- 0010011000010010  not	r2, r2
  691=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  692=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  693=>x"D221",	-- 1101001000100001  sw	r1, r4
  694=>x"C0A1",	-- 1100000010100001  li	r1, 20
  695=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  696=>x"D03A",	-- 1101000000111010  lw	r2, r7
  697=>x"043F",	-- 0000010000111111  inc	r7, r7
  698=>x"0412",	-- 0000010000010010  inc	r2, r2
  699=>x"061B",	-- 0000011000011011  dec	r3, r3
  700=>x"E398",	-- 1110001110011000  baeq	r3, r6
  701=>x"B683",	-- 1011011010000011  bri	-, put_sprite_8.loop0
  702=>x"D010",	-- 1101000000010000  lw	r0, r2
  703=>x"063F",	-- 0000011000111111  dec	r7, r7
  704=>x"D23A",	-- 1101001000111010  sw	r2, r7
  705=>x"063F",	-- 0000011000111111  dec	r7, r7
  706=>x"D23B",	-- 1101001000111011  sw	r3, r7
  707=>x"C802",	-- 1100100000000010  li	r2, 0x100
  708=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  709=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  710=>x"2080",	-- 0010000010000000  and	r0, r0, r2
  711=>x"D021",	-- 1101000000100001  lw	r1, r4
  712=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
  713=>x"261B",	-- 0010011000011011  not	r3, r3
  714=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  715=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
  716=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  717=>x"D221",	-- 1101001000100001  sw	r1, r4
  718=>x"0424",	-- 0000010000100100  inc	r4, r4
  719=>x"D021",	-- 1101000000100001  lw	r1, r4
  720=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  721=>x"261B",	-- 0010011000011011  not	r3, r3
  722=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  723=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
  724=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  725=>x"D221",	-- 1101001000100001  sw	r1, r4
  726=>x"C099",	-- 1100000010011001  li	r1, 19
  727=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  728=>x"D03B",	-- 1101000000111011  lw	r3, r7
  729=>x"043F",	-- 0000010000111111  inc	r7, r7
  730=>x"D03A",	-- 1101000000111010  lw	r2, r7
  731=>x"043F",	-- 0000010000111111  inc	r7, r7
  732=>x"061B",	-- 0000011000011011  dec	r3, r3
  733=>x"E398",	-- 1110001110011000  baeq	r3, r6
  734=>x"D010",	-- 1101000000010000  lw	r0, r2
  735=>x"4E00",	-- 0100111000000000  shl	r0, r0, 7
  736=>x"063F",	-- 0000011000111111  dec	r7, r7
  737=>x"D23A",	-- 1101001000111010  sw	r2, r7
  738=>x"063F",	-- 0000011000111111  dec	r7, r7
  739=>x"D23B",	-- 1101001000111011  sw	r3, r7
  740=>x"C802",	-- 1100100000000010  li	r2, 0x100
  741=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  742=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  743=>x"2080",	-- 0010000010000000  and	r0, r0, r2
  744=>x"D021",	-- 1101000000100001  lw	r1, r4
  745=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
  746=>x"261B",	-- 0010011000011011  not	r3, r3
  747=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  748=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
  749=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  750=>x"D221",	-- 1101001000100001  sw	r1, r4
  751=>x"0424",	-- 0000010000100100  inc	r4, r4
  752=>x"D021",	-- 1101000000100001  lw	r1, r4
  753=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  754=>x"261B",	-- 0010011000011011  not	r3, r3
  755=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  756=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
  757=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  758=>x"D221",	-- 1101001000100001  sw	r1, r4
  759=>x"C099",	-- 1100000010011001  li	r1, 19
  760=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  761=>x"D03B",	-- 1101000000111011  lw	r3, r7
  762=>x"043F",	-- 0000010000111111  inc	r7, r7
  763=>x"D03A",	-- 1101000000111010  lw	r2, r7
  764=>x"043F",	-- 0000010000111111  inc	r7, r7
  765=>x"0412",	-- 0000010000010010  inc	r2, r2
  766=>x"061B",	-- 0000011000011011  dec	r3, r3
  767=>x"E398",	-- 1110001110011000  baeq	r3, r6
  768=>x"AF83",	-- 1010111110000011  bri	-, put_sprite_8.loop1
    others => x"0000"
    );
begin
  process(CLK)
  begin
    if (CLK'event AND CLK='1') then
      D <= m(to_integer(unsigned(AD)));
    end if;
  end process;
end Behavioral;
