----------------------------------------------------------------------------------
--
-- File retrieved, on 07/02/2010, from :
-- http://sebastien-viardot.imag.fr/Enseignements/Archi1A2s/sources/ROMPROG.vhd
--
-- Slightly altered to get rid of vendor-specific packages and adjust formatting
-- Now auto-filled by asrom script
--
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROMPROG is
  Port ( AD : in  STD_LOGIC_VECTOR (12 downto 0);
         D : out  STD_LOGIC_VECTOR (15 downto 0);
         CLK : in STD_LOGIC);
end ROMPROG;

architecture Behavioral of ROMPROG is
  constant low_address: natural := 0;
  constant high_address: natural := 8192;
  subtype octet is std_logic_vector( 15 downto 0 );
  type zone_memoire is
    array (natural range low_address to high_address-1) of octet;
  constant m: zone_memoire:= (
    0=>x"FFF7",	-- 1111111111110111  liw	r7, IRQ_mask
    1=>x"2000",	-- 0010000000000000  
    2=>x"F8C0",	-- 1111100011000000  bai	-, os_init
    3=>x"0100",	-- 0000000100000000  
   16=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_ack
   17=>x"2002",	-- 0010000000000010  
   18=>x"D001",	-- 1101000000000001  lw	r1, r0
   19=>x"F54A",	-- 1111010101001010  bspl	r2, r1, 5
   20=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_error
   21=>x"0050",	-- 0000000001010000  
   22=>x"F4CA",	-- 1111010011001010  bspl	r2, r1, 3
   23=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_kbd
   24=>x"0060",	-- 0000000001100000  
   25=>x"F40A",	-- 1111010000001010  bspl	r2, r1, 0
   26=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_tmr
   27=>x"0040",	-- 0000000001000000  
   28=>x"D201",	-- 1101001000000001  sw	r1, r0
   29=>x"FFFE",	-- 1111111111111110  reti
   64=>x"263F",	-- 0010011000111111  not r7, r7
   65=>x"D7C0",	-- 1101011111000000  out	r7
   66=>x"E383",	-- 1110001110000011  ba	-, r6
   80=>x"25FF",	-- 0010010111111111  xor	r7, r7, r7
   81=>x"D7C0",	-- 1101011111000000  out	r7
   82=>x"E383",	-- 1110001110000011  ba	-, r6
   96=>x"FFF2",	-- 1111111111110010  liw	r2, PS2_rx
   97=>x"2004",	-- 0010000000000100  
   98=>x"D012",	-- 1101000000010010  lw	r2, r2
   99=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map + 8
  100=>x"16C8",	-- 0001011011001000  
  101=>x"D01B",	-- 1101000000011011  lw	r3, r3
  102=>x"1EBF",	-- 0001111010111111  mixll	r7, r7, r2
  103=>x"C784",	-- 1100011110000100  li	r4, 0xF0
  104=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  105=>x"8C60",	-- 1000110001100000  brieq	r4, int_kbd.release
  106=>x"C704",	-- 1100011100000100  li	r4, 0xE0
  107=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  108=>x"8A20",	-- 1000101000100000  brieq	r4, int_kbd.extended
  109=>x"FFF5",	-- 1111111111110101  liw	r5, rand_seed
  110=>x"16C8",	-- 0001011011001000  
  111=>x"D02C",	-- 1101000000101100  lw	r4, r5
  112=>x"24A4",	-- 0010010010100100  xor	r4, r4, r2
  113=>x"D22C",	-- 1101001000101100  sw	r4, r5
  114=>x"FFF5",	-- 1111111111110101  liw	r5, paper_keys - 1
  115=>x"16CF",	-- 0001011011001111  
  116=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  117=>x"80E0",	-- 1000000011100000  brieq	r4, $+3
  118=>x"FFF5",	-- 1111111111110101  liw	r5, paper_keys + 11 - 1
  119=>x"16DA",	-- 0001011011011010  
  120=>x"042D",	-- 0000010000101101  inc	r5, r5
  121=>x"D02C",	-- 1101000000101100  lw	r4, r5
  122=>x"8560",	-- 1000010101100000  brieq	r4, scan_code_mismatch
  123=>x"6E24",	-- 0110111000100100  shr	r4, r4, 7
  124=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  125=>x"BEE4",	-- 1011111011100100  brine	r4, scan_code_loop
  126=>x"D02A",	-- 1101000000101010  lw	r2, r5
  127=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  128=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  129=>x"741B",	-- 0111010000011011  shr	r3, r3, 10
  130=>x"C00D",	-- 1100000000001101  li	r5, 1
  131=>x"0612",	-- 0000011000010010  dec	r2, r2
  132=>x"3AAA",	-- 0011101010101010  rrl	r2, r5, r2
  133=>x"FFF5",	-- 1111111111110101  liw	r5, key_press_map
  134=>x"16C0",	-- 0001011011000000  
  135=>x"08ED",	-- 0000100011101101  add	r5, r5, r3
  136=>x"D02B",	-- 1101000000101011  lw	r3, r5
  137=>x"80E4",	-- 1000000011100100  brine	r4, scan_code_release
  138=>x"229B",	-- 0010001010011011  or	r3, r3, r2
  139=>x"80C3",	-- 1000000011000011  bri	-, scan_code_notify
  140=>x"2612",	-- 0010011000010010  not	r2, r2
  141=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  142=>x"D22B",	-- 1101001000101011  sw	r3, r5
  143=>x"C003",	-- 1100000000000011  li	r3, 0
  144=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  145=>x"16C8",	-- 0001011011001000  
  146=>x"D223",	-- 1101001000100011  sw	r3, r4
  147=>x"E383",	-- 1110001110000011  ba	-, r6
  148=>x"C014",	-- 1100000000010100  li	r4, 2
  149=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  150=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  151=>x"16C8",	-- 0001011011001000  
  152=>x"D223",	-- 1101001000100011  sw	r3, r4
  153=>x"E383",	-- 1110001110000011  ba	-, r6
  154=>x"C00C",	-- 1100000000001100  li	r4, 1
  155=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  156=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  157=>x"16C8",	-- 0001011011001000  
  158=>x"D223",	-- 1101001000100011  sw	r3, r4
  159=>x"E383",	-- 1110001110000011  ba	-, r6
  256=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_mask
  257=>x"2000",	-- 0010000000000000  
  258=>x"C0C9",	-- 1100000011001001  li	r1, 0x19
  259=>x"D201",	-- 1101001000000001  sw	r1, r0
  260=>x"0400",	-- 0000010000000000  inc	r0, r0
  261=>x"CFF9",	-- 1100111111111001  li	r1, -1
  262=>x"D201",	-- 1101001000000001  sw	r1, r0
  263=>x"C03A",	-- 1100000000111010  li	r2, 7
  264=>x"0880",	-- 0000100010000000  add	r0, r0, r2
  265=>x"C0EA",	-- 1100000011101010  li	r2, 0x1D
  266=>x"D202",	-- 1101001000000010  sw	r2, r0
  267=>x"0400",	-- 0000010000000000  inc	r0, r0
  268=>x"C07A",	-- 1100000001111010  li	r2, 15
  269=>x"D202",	-- 1101001000000010  sw	r2, r0
  270=>x"0400",	-- 0000010000000000  inc	r0, r0
  271=>x"C0DA",	-- 1100000011011010  li	r2, 0x1B
  272=>x"D202",	-- 1101001000000010  sw	r2, r0
  273=>x"0400",	-- 0000010000000000  inc	r0, r0
  274=>x"FFF2",	-- 1111111111110010  liw	r2, 817
  275=>x"0331",	-- 0000001100110001  
  276=>x"D202",	-- 1101001000000010  sw	r2, r0
  277=>x"FFF0",	-- 1111111111110000  liw	r0, key_press_map
  278=>x"16C0",	-- 0001011011000000  
  279=>x"C001",	-- 1100000000000001  li	r1, 0
  280=>x"C042",	-- 1100000001000010  li	r2, 8
  281=>x"D201",	-- 1101001000000001  sw	r1, r0
  282=>x"0400",	-- 0000010000000000  inc	r0, r0
  283=>x"0612",	-- 0000011000010010  dec	r2, r2
  284=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  285=>x"8083",	-- 1000000010000011  bri	-, PaperGameStart
  286=>x"8003",	-- 1000000000000011  bri	-, PaperMenuLoop
  287=>x"FFF0",	-- 1111111111110000  liw	r0, paper_dir
  288=>x"179C",	-- 0001011110011100  
  289=>x"C001",	-- 1100000000000001  li	r1, 0
  290=>x"D201",	-- 1101001000000001  sw	r1, r0
  291=>x"0400",	-- 0000010000000000  inc	r0, r0
  292=>x"FFF1",	-- 1111111111110001  liw	r1, 152 * 8
  293=>x"04C0",	-- 0000010011000000  
  294=>x"D201",	-- 1101001000000001  sw	r1, r0
  295=>x"0400",	-- 0000010000000000  inc	r0, r0
  296=>x"C001",	-- 1100000000000001  li	r1, 0
  297=>x"D201",	-- 1101001000000001  sw	r1, r0
  298=>x"0400",	-- 0000010000000000  inc	r0, r0
  299=>x"FFF1",	-- 1111111111110001  liw	r1, 128 * 8
  300=>x"0400",	-- 0000010000000000  
  301=>x"D201",	-- 1101001000000001  sw	r1, r0
  302=>x"0400",	-- 0000010000000000  inc	r0, r0
  303=>x"C001",	-- 1100000000000001  li	r1, 0
  304=>x"D201",	-- 1101001000000001  sw	r1, r0
  305=>x"0400",	-- 0000010000000000  inc	r0, r0
  306=>x"C069",	-- 1100000001101001  li	r1, 13
  307=>x"D201",	-- 1101001000000001  sw	r1, r0
  308=>x"0400",	-- 0000010000000000  inc	r0, r0
  309=>x"C011",	-- 1100000000010001  li	r1, 2
  310=>x"D201",	-- 1101001000000001  sw	r1, r0
  311=>x"0400",	-- 0000010000000000  inc	r0, r0
  312=>x"FFF0",	-- 1111111111110000  liw	r0, paper_tilemap
  313=>x"17B0",	-- 0001011110110000  
  314=>x"C001",	-- 1100000000000001  li	r1, 0
  315=>x"C0C2",	-- 1100000011000010  li	r2, 6*4
  316=>x"D201",	-- 1101001000000001  sw	r1, r0
  317=>x"0400",	-- 0000010000000000  inc	r0, r0
  318=>x"0612",	-- 0000011000010010  dec	r2, r2
  319=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  320=>x"C000",	-- 1100000000000000  li	r0, 0
  321=>x"CFF9",	-- 1100111111111001  li	r1, -1
  322=>x"C0A2",	-- 1100000010100010  li	r2, 20
  323=>x"D201",	-- 1101001000000001  sw	r1, r0
  324=>x"0400",	-- 0000010000000000  inc	r0, r0
  325=>x"0612",	-- 0000011000010010  dec	r2, r2
  326=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  327=>x"C001",	-- 1100000000000001  li	r1, 0
  328=>x"FFF2",	-- 1111111111110010  liw	r2, 18*20
  329=>x"0168",	-- 0000000101101000  
  330=>x"D201",	-- 1101001000000001  sw	r1, r0
  331=>x"0400",	-- 0000010000000000  inc	r0, r0
  332=>x"0612",	-- 0000011000010010  dec	r2, r2
  333=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  334=>x"CFF9",	-- 1100111111111001  li	r1, -1
  335=>x"C0A2",	-- 1100000010100010  li	r2, 20
  336=>x"D201",	-- 1101001000000001  sw	r1, r0
  337=>x"0400",	-- 0000010000000000  inc	r0, r0
  338=>x"0612",	-- 0000011000010010  dec	r2, r2
  339=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  340=>x"C020",	-- 1100000000100000  li	r0, 4
  341=>x"C029",	-- 1100000000101001  li	r1, 5
  342=>x"FFF2",	-- 1111111111110010  liw	r2, paper_title
  343=>x"17A4",	-- 0001011110100100  
  344=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  345=>x"02A9",	-- 0000001010101001  
  346=>x"C090",	-- 1100000010010000  li	r0, 18
  347=>x"C029",	-- 1100000000101001  li	r1, 5
  348=>x"FFF2",	-- 1111111111110010  liw	r2, paper_score
  349=>x"16C9",	-- 0001011011001001  
  350=>x"D012",	-- 1101000000010010  lw	r2, r2
  351=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum
  352=>x"02D8",	-- 0000001011011000  
  353=>x"C778",	-- 1100011101111000  li	r0, 239
  354=>x"C009",	-- 1100000000001001  li	r1, 1
  355=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud
  356=>x"1780",	-- 0001011110000000  
  357=>x"C043",	-- 1100000001000011  li	r3, 8
  358=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  359=>x"03B1",	-- 0000001110110001  
  360=>x"C0F8",	-- 1100000011111000  li	r0, 31
  361=>x"C009",	-- 1100000000001001  li	r1, 1
  362=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  363=>x"17A0",	-- 0001011110100000  
  364=>x"D012",	-- 1101000000010010  lw	r2, r2
  365=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum
  366=>x"02D8",	-- 0000001011011000  
  367=>x"C120",	-- 1100000100100000  li	r0, 36
  368=>x"C009",	-- 1100000000001001  li	r1, 1
  369=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  370=>x"17AA",	-- 0001011110101010  
  371=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  372=>x"02A9",	-- 0000001010101001  
  373=>x"C778",	-- 1100011101111000  li	r0, 239
  374=>x"C051",	-- 1100000001010001  li	r1, 10
  375=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud + 8
  376=>x"1788",	-- 0001011110001000  
  377=>x"C043",	-- 1100000001000011  li	r3, 8
  378=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  379=>x"03B1",	-- 0000001110110001  
  380=>x"C0F8",	-- 1100000011111000  li	r0, 31
  381=>x"C051",	-- 1100000001010001  li	r1, 10
  382=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed + 1
  383=>x"17A1",	-- 0001011110100001  
  384=>x"D012",	-- 1101000000010010  lw	r2, r2
  385=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum
  386=>x"02D8",	-- 0000001011011000  
  387=>x"C120",	-- 1100000100100000  li	r0, 36
  388=>x"C051",	-- 1100000001010001  li	r1, 10
  389=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  390=>x"17AA",	-- 0001011110101010  
  391=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  392=>x"02A9",	-- 0000001010101001  
  393=>x"FFF0",	-- 1111111111110000  liw	r0, 20*20
  394=>x"0190",	-- 0000000110010000  
  395=>x"C001",	-- 1100000000000001  li	r1, 0
  396=>x"FFF2",	-- 1111111111110010  liw	r2, 220*20
  397=>x"1130",	-- 0001000100110000  
  398=>x"D201",	-- 1101001000000001  sw	r1, r0
  399=>x"0400",	-- 0000010000000000  inc	r0, r0
  400=>x"0612",	-- 0000011000010010  dec	r2, r2
  401=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  402=>x"FFF5",	-- 1111111111110101  liw	r5, paper_tilemap
  403=>x"17B0",	-- 0001011110110000  
  404=>x"D02C",	-- 1101000000101100  lw	r4, r5
  405=>x"042D",	-- 0000010000101101  inc	r5, r5
  406=>x"8960",	-- 1000100101100000  brieq	r4, PaperGameTileSkip
  407=>x"063F",	-- 0000011000111111  dec	r7, r7
  408=>x"D23D",	-- 1101001000111101  sw	r5, r7
  409=>x"FFF3",	-- 1111111111110011  liw	r3, paper_tilemap
  410=>x"17B0",	-- 0001011110110000  
  411=>x"0AEB",	-- 0000101011101011  sub	r3, r5, r3
  412=>x"6E20",	-- 0110111000100000  shr	r0, r4, 7
  413=>x"6219",	-- 0110001000011001  shr	r1, r3, 1
  414=>x"4809",	-- 0100100000001001  shl	r1, r1, 4
  415=>x"C19A",	-- 1100000110011010  li	r2, 51
  416=>x"0889",	-- 0000100010001001  add	r1, r1, r2
  417=>x"FFF2",	-- 1111111111110010  liw	r2, paper_pos + 1
  418=>x"179E",	-- 0001011110011110  
  419=>x"D012",	-- 1101000000010010  lw	r2, r2
  420=>x"6412",	-- 0110010000010010  shr	r2, r2, 2
  421=>x"C0FB",	-- 1100000011111011  li	r3, 31
  422=>x"20D2",	-- 0010000011010010  and	r2, r2, r3
  423=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  424=>x"4E24",	-- 0100111000100100  shl	r4, r4, 7
  425=>x"6E24",	-- 0110111000100100  shr	r4, r4, 7
  426=>x"C00B",	-- 1100000000001011  li	r3, 1
  427=>x"FB06",	-- 1111101100000110  bailne	r0, r6, put_tile
  428=>x"0279",	-- 0000001001111001  
  429=>x"81E0",	-- 1000000111100000  brieq	r4, PaperGameSegmentSkip
  431=>x"C013",	-- 1100000000010011  li	r3, 2
  432=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_tile
  433=>x"0279",	-- 0000001001111001  
  434=>x"0624",	-- 0000011000100100  dec	r4, r4
  435=>x"BF64",	-- 1011111101100100  brine	r4, PaperGameSegmentLoop
  436=>x"C003",	-- 1100000000000011  li	r3, 0
  437=>x"C144",	-- 1100000101000100  li	r4, 40
  438=>x"0B04",	-- 0000101100000100  sub	r4, r0, r4
  439=>x"FB66",	-- 1111101101100110  baillt	r4, r6, put_tile
  440=>x"0279",	-- 0000001001111001  
  441=>x"D03D",	-- 1101000000111101  lw	r5, r7
  442=>x"043F",	-- 0000010000111111  inc	r7, r7
  443=>x"FFF4",	-- 1111111111110100  liw r4, paper_tilemap + 24
  444=>x"17C8",	-- 0001011111001000  
  445=>x"0B2C",	-- 0000101100101100  sub	r4, r5, r4
  446=>x"B5A5",	-- 1011010110100101  brilt	r4, PaperGameTileLoop
  447=>x"FFF3",	-- 1111111111110011  liw	r3, paper_speed
  448=>x"17A0",	-- 0001011110100000  
  449=>x"D01B",	-- 1101000000011011  lw	r3, r3
  450=>x"CF04",	-- 1100111100000100  li	r4, 0x1E0
  451=>x"211C",	-- 0010000100011100  and	r4, r3, r4
  452=>x"FFF3",	-- 1111111111110011  liw	r3, paper_pos
  453=>x"179D",	-- 0001011110011101  
  454=>x"D018",	-- 1101000000011000  lw	r0, r3
  455=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  456=>x"FFF2",	-- 1111111111110010  liw	r2, paper_sprites
  457=>x"1720",	-- 0001011100100000  
  458=>x"0912",	-- 0000100100010010  add	r2, r2, r4
  459=>x"C161",	-- 1100000101100001  li	r1, 44
  460=>x"C083",	-- 1100000010000011  li	r3, 16
  461=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_16_masked
  462=>x"0349",	-- 0000001101001001  
  463=>x"912C",	-- 1001000100101100  brine	r5, PaperGameFail
  465=>x"C028",	-- 1100000000101000  li	r0, 5
  466=>x"C001",	-- 1100000000000001  li	r1, 0
  467=>x"8043",	-- 1000000001000011  bri	-, $+1
  468=>x"0609",	-- 0000011000001001  dec	r1, r1
  469=>x"BF8C",	-- 1011111110001100  brine	r1, $-2
  470=>x"0600",	-- 0000011000000000  dec	r0, r0
  471=>x"BEC4",	-- 1011111011000100  brine	r0, $-5
  472=>x"FFF2",	-- 1111111111110010  liw	r2, paper_pos
  473=>x"179D",	-- 0001011110011101  
  474=>x"FFF3",	-- 1111111111110011  liw	r3, paper_speed
  475=>x"17A0",	-- 0001011110100000  
  476=>x"D010",	-- 1101000000010000  lw	r0, r2
  477=>x"D019",	-- 1101000000011001  lw	r1, r3
  478=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  479=>x"8D05",	-- 1000110100000101  brilt	r0, PaperGameFail
  480=>x"FFF4",	-- 1111111111110100  liw	r4, 304*8
  481=>x"0980",	-- 0000100110000000  
  482=>x"0B04",	-- 0000101100000100  sub	r4, r0, r4
  483=>x"8C21",	-- 1000110000100001  brige	r4, PaperGameFail
  484=>x"D210",	-- 1101001000010000  sw	r0, r2
  485=>x"F7CD",	-- 1111011111001101  bspl	r5, r1, 15
  486=>x"80A8",	-- 1000000010101000  brieq	r5, $+2
  487=>x"1409",	-- 0001010000001001  nega	r1, r1
  488=>x"660D",	-- 0110011000001101  shr	r5, r1, 3
  489=>x"0412",	-- 0000010000010010  inc	r2, r2
  490=>x"041B",	-- 0000010000011011  inc	r3, r3
  491=>x"D010",	-- 1101000000010000  lw	r0, r2
  492=>x"D019",	-- 1101000000011001  lw	r1, r3
  493=>x"C7FC",	-- 1100011111111100  li	r4, 0xFF
  494=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  495=>x"0B40",	-- 0000101101000000  sub	r0, r0, r5
  496=>x"2101",	-- 0010000100000001  and	r1, r0, r4
  497=>x"D211",	-- 1101001000010001  sw	r1, r2
  498=>x"2624",	-- 0010011000100100  not	r4, r4
  499=>x"2100",	-- 0010000100000000  and	r0, r0, r4
  500=>x"FB06",	-- 1111101100000110  bailne	r0, r6, PaperMapScroll
  501=>x"0221",	-- 0000001000100001  
  502=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  503=>x"16C0",	-- 0001011011000000  
  504=>x"D01B",	-- 1101000000011011  lw	r3, r3
  505=>x"F818",	-- 1111100000011000  baieq	r3, PaperGameRedraw
  506=>x"0140",	-- 0000000101000000  
  507=>x"F7DC",	-- 1111011111011100  bspl	r4, r3, 15
  508=>x"8924",	-- 1000100100100100  brine	r4, PaperGameQuit
  509=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  510=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveUp
  511=>x"F49C",	-- 1111010010011100  bspl	r4, r3, 2
  512=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveDOWN
  513=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  514=>x"81E0",	-- 1000000111100000  brieq	r4, PaperNoMoveLEFT
  515=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  516=>x"17A0",	-- 0001011110100000  
  517=>x"D010",	-- 1101000000010000  lw	r0, r2
  518=>x"C02C",	-- 1100000000101100  li	r4, 5
  519=>x"0B00",	-- 0000101100000000  sub	r0, r0, r4
  520=>x"D210",	-- 1101001000010000  sw	r0, r2
  521=>x"F4DC",	-- 1111010011011100  bspl	r4, r3, 3
  522=>x"81E0",	-- 1000000111100000  brieq	r4, PaperNoMoveRIGHT
  523=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  524=>x"17A0",	-- 0001011110100000  
  525=>x"D010",	-- 1101000000010000  lw	r0, r2
  526=>x"C02C",	-- 1100000000101100  li	r4, 5
  527=>x"0900",	-- 0000100100000000  add	r0, r0, r4
  528=>x"D210",	-- 1101001000010000  sw	r0, r2
  529=>x"F8C0",	-- 1111100011000000  bai	-, PaperGameRedraw
  530=>x"0140",	-- 0000000101000000  
  531=>x"C000",	-- 1100000000000000  li	r0, 0
  532=>x"FFF2",	-- 1111111111110010  liw	r2, 240*20
  533=>x"12C0",	-- 0001001011000000  
  534=>x"D001",	-- 1101000000000001  lw	r1, r0
  535=>x"2609",	-- 0010011000001001  not	r1, r1
  536=>x"D201",	-- 1101001000000001  sw	r1, r0
  537=>x"0400",	-- 0000010000000000  inc	r0, r0
  538=>x"0612",	-- 0000011000010010  dec	r2, r2
  539=>x"BED4",	-- 1011111011010100  brine	r2, $-5
  540=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  541=>x"16C0",	-- 0001011011000000  
  542=>x"D01A",	-- 1101000000011010  lw	r2, r3
  543=>x"BFD0",	-- 1011111111010000  brieq	r2, $-1
  544=>x"FFFF",	-- 1111111111111111  reset
  545=>x"FFF0",	-- 1111111111110000  liw	r0, paper_tilemap
  546=>x"17B0",	-- 0001011110110000  
  547=>x"C021",	-- 1100000000100001  li	r1, 4
  548=>x"0841",	-- 0000100001000001  add	r1, r0, r1
  549=>x"C0A2",	-- 1100000010100010  li	r2, 5*4
  550=>x"D00B",	-- 1101000000001011  lw	r3, r1
  551=>x"D203",	-- 1101001000000011  sw	r3, r0
  552=>x"0400",	-- 0000010000000000  inc	r0, r0
  553=>x"0409",	-- 0000010000001001  inc	r1, r1
  554=>x"0612",	-- 0000011000010010  dec	r2, r2
  555=>x"BED4",	-- 1011111011010100  brine	r2, PaperGameScrollLoop
  556=>x"063F",	-- 0000011000111111  dec	r7, r7
  557=>x"D23E",	-- 1101001000111110  sw	r6, r7
  558=>x"FAC6",	-- 1111101011000110  bail	-, r6, rand16
  559=>x"0267",	-- 0000001001100111  
  560=>x"C02A",	-- 1100000000101010  li	r2, 0x05
  561=>x"208B",	-- 0010000010001011  and	r3, r1, r2
  562=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  563=>x"208C",	-- 0010000010001100  and	r4, r1, r2
  564=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  565=>x"1F19",	-- 0001111100011001  mixll	r1, r3, r4
  566=>x"D201",	-- 1101001000000001  sw	r1, r0
  567=>x"0400",	-- 0000010000000000  inc	r0, r0
  568=>x"C03A",	-- 1100000000111010  li	r2, 0x07
  569=>x"091C",	-- 0000100100011100  add r4, r3, r4
  570=>x"208B",	-- 0010000010001011  and	r3, r1, r2
  571=>x"091C",	-- 0000100100011100  add r4, r3, r4
  572=>x"C01B",	-- 1100000000011011  li	r3, 3
  573=>x"08E4",	-- 0000100011100100  add	r4, r4, r3
  574=>x"6209",	-- 0110001000001001  shr	r1, r1, 1
  575=>x"208B",	-- 0010000010001011  and	r3, r1, r2
  576=>x"091B",	-- 0000100100011011  add r3, r3, r4
  577=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  578=>x"208C",	-- 0010000010001100  and	r4, r1, r2
  579=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  580=>x"1F19",	-- 0001111100011001  mixll	r1, r3, r4
  581=>x"D201",	-- 1101001000000001  sw	r1, r0
  582=>x"0400",	-- 0000010000000000  inc	r0, r0
  583=>x"C02A",	-- 1100000000101010  li	r2, 0x05
  584=>x"091C",	-- 0000100100011100  add r4, r3, r4
  585=>x"208B",	-- 0010000010001011  and	r3, r1, r2
  586=>x"091C",	-- 0000100100011100  add r4, r3, r4
  587=>x"C01B",	-- 1100000000011011  li	r3, 3
  588=>x"08E4",	-- 0000100011100100  add	r4, r4, r3
  589=>x"6209",	-- 0110001000001001  shr	r1, r1, 1
  590=>x"208B",	-- 0010000010001011  and	r3, r1, r2
  591=>x"091B",	-- 0000100100011011  add r3, r3, r4
  592=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  593=>x"208C",	-- 0010000010001100  and	r4, r1, r2
  594=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  595=>x"1F19",	-- 0001111100011001  mixll	r1, r3, r4
  596=>x"D201",	-- 1101001000000001  sw	r1, r0
  597=>x"0400",	-- 0000010000000000  inc	r0, r0
  598=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed + 1
  599=>x"17A1",	-- 0001011110100001  
  600=>x"D011",	-- 1101000000010001  lw	r1, r2
  601=>x"0409",	-- 0000010000001001  inc	r1, r1
  602=>x"D211",	-- 1101001000010001  sw	r1, r2
  603=>x"FFF2",	-- 1111111111110010  liw	r2, paper_score
  604=>x"16C9",	-- 0001011011001001  
  605=>x"D011",	-- 1101000000010001  lw	r1, r2
  606=>x"0409",	-- 0000010000001001  inc	r1, r1
  607=>x"D211",	-- 1101001000010001  sw	r1, r2
  608=>x"D03E",	-- 1101000000111110  lw	r6, r7
  609=>x"043F",	-- 0000010000111111  inc	r7, r7
  610=>x"E383",	-- 1110001110000011  ba	-, r6
  611=>x"FFF2",	-- 1111111111110010  liw	r2, rand_seed
  612=>x"16C8",	-- 0001011011001000  
  613=>x"D210",	-- 1101001000010000  sw	r0, r2
  614=>x"E383",	-- 1110001110000011  ba	-, r6
  615=>x"FFF2",	-- 1111111111110010  liw	r2, rand_seed
  616=>x"16C8",	-- 0001011011001000  
  617=>x"D013",	-- 1101000000010011  lw	r3, r2
  618=>x"C7EC",	-- 1100011111101100  li	r4, 253
  619=>x"1F19",	-- 0001111100011001  mixll	r1, r3, r4
  620=>x"18E4",	-- 0001100011100100  mixhh	r4, r4, r3
  621=>x"C002",	-- 1100000000000010  li	r2, 0
  622=>x"0AC9",	-- 0000101011001001  sub	r1, r1, r3
  623=>x"0EA4",	-- 0000111010100100  sbc	r4, r4, r2
  624=>x"0EC9",	-- 0000111011001001  sbc	r1, r1, r3
  625=>x"0EA4",	-- 0000111010100100  sbc	r4, r4, r2
  626=>x"1B13",	-- 0001101100010011  mixhl	r3, r2, r4
  627=>x"0EC9",	-- 0000111011001001  sbc	r1, r1, r3
  628=>x"0C89",	-- 0000110010001001  adc	r1, r1, r2
  629=>x"FFF2",	-- 1111111111110010  liw	r2, rand_seed
  630=>x"16C8",	-- 0001011011001000  
  631=>x"D211",	-- 1101001000010001  sw	r1, r2
  632=>x"E383",	-- 1110001110000011  ba	-, r6
  633=>x"063F",	-- 0000011000111111  dec	r7, r7
  634=>x"D238",	-- 1101001000111000  sw	r0, r7
  635=>x"063F",	-- 0000011000111111  dec	r7, r7
  636=>x"D239",	-- 1101001000111001  sw	r1, r7
  637=>x"063F",	-- 0000011000111111  dec	r7, r7
  638=>x"D23A",	-- 1101001000111010  sw	r2, r7
  639=>x"063F",	-- 0000011000111111  dec	r7, r7
  640=>x"D23B",	-- 1101001000111011  sw	r3, r7
  641=>x"063F",	-- 0000011000111111  dec	r7, r7
  642=>x"D23C",	-- 1101001000111100  sw	r4, r7
  643=>x"063F",	-- 0000011000111111  dec	r7, r7
  644=>x"D23D",	-- 1101001000111101  sw	r5, r7
  645=>x"063F",	-- 0000011000111111  dec	r7, r7
  646=>x"D23E",	-- 1101001000111110  sw	r6, r7
  647=>x"FFF2",	-- 1111111111110010  liw	r2, paper_tiles
  648=>x"1790",	-- 0001011110010000  
  649=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  650=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  651=>x"C043",	-- 1100000001000011  li	r3, 8
  652=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  653=>x"038B",	-- 0000001110001011  
  654=>x"D03E",	-- 1101000000111110  lw	r6, r7
  655=>x"043F",	-- 0000010000111111  inc	r7, r7
  656=>x"D03D",	-- 1101000000111101  lw	r5, r7
  657=>x"043F",	-- 0000010000111111  inc	r7, r7
  658=>x"D03C",	-- 1101000000111100  lw	r4, r7
  659=>x"043F",	-- 0000010000111111  inc	r7, r7
  660=>x"D03B",	-- 1101000000111011  lw	r3, r7
  661=>x"043F",	-- 0000010000111111  inc	r7, r7
  662=>x"D03A",	-- 1101000000111010  lw	r2, r7
  663=>x"043F",	-- 0000010000111111  inc	r7, r7
  664=>x"D039",	-- 1101000000111001  lw	r1, r7
  665=>x"043F",	-- 0000010000111111  inc	r7, r7
  666=>x"D038",	-- 1101000000111000  lw	r0, r7
  667=>x"043F",	-- 0000010000111111  inc	r7, r7
  668=>x"0400",	-- 0000010000000000  inc	r0, r0
  669=>x"E383",	-- 1110001110000011  ba	-, r6
  670=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  671=>x"C084",	-- 1100000010000100  li	r4, 16
  672=>x"0800",	-- 0000100000000000  add	r0, r0, r0
  673=>x"0C49",	-- 0000110001001001  adc	r1, r1, r1
  674=>x"0A8B",	-- 0000101010001011  sub	r3, r1, r2
  675=>x"80DD",	-- 1000000011011101  brilt	r3, div_16_16.skip
  676=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  677=>x"0400",	-- 0000010000000000  inc	r0, r0
  678=>x"0624",	-- 0000011000100100  dec	r4, r4
  679=>x"BE64",	-- 1011111001100100  brine	r4, div_16_16.loop
  680=>x"E383",	-- 1110001110000011  ba	-, r6
  681=>x"063F",	-- 0000011000111111  dec	r7, r7
  682=>x"D23E",	-- 1101001000111110  sw	r6, r7
  683=>x"D013",	-- 1101000000010011  lw	r3, r2
  684=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  685=>x"84D8",	-- 1000010011011000  brieq	r3, puts.end
  686=>x"063F",	-- 0000011000111111  dec	r7, r7
  687=>x"D23A",	-- 1101001000111010  sw	r2, r7
  688=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  689=>x"02C3",	-- 0000001011000011  
  690=>x"D03A",	-- 1101000000111010  lw	r2, r7
  691=>x"043F",	-- 0000010000111111  inc	r7, r7
  692=>x"D013",	-- 1101000000010011  lw	r3, r2
  693=>x"4E1B",	-- 0100111000011011  shl	r3, r3, 7
  694=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  695=>x"8258",	-- 1000001001011000  brieq	r3, puts.end
  696=>x"063F",	-- 0000011000111111  dec	r7, r7
  697=>x"D23A",	-- 1101001000111010  sw	r2, r7
  698=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  699=>x"02C3",	-- 0000001011000011  
  700=>x"D03A",	-- 1101000000111010  lw	r2, r7
  701=>x"043F",	-- 0000010000111111  inc	r7, r7
  702=>x"0412",	-- 0000010000010010  inc	r2, r2
  703=>x"BB03",	-- 1011101100000011  bri	-, puts.loop
  704=>x"D03E",	-- 1101000000111110  lw	r6, r7
  705=>x"043F",	-- 0000010000111111  inc	r7, r7
  706=>x"E383",	-- 1110001110000011  ba	-, r6
  707=>x"063F",	-- 0000011000111111  dec	r7, r7
  708=>x"D23E",	-- 1101001000111110  sw	r6, r7
  709=>x"063F",	-- 0000011000111111  dec	r7, r7
  710=>x"D238",	-- 1101001000111000  sw	r0, r7
  711=>x"063F",	-- 0000011000111111  dec	r7, r7
  712=>x"D239",	-- 1101001000111001  sw	r1, r7
  713=>x"FFF2",	-- 1111111111110010  liw	r2, font_map
  714=>x"12C0",	-- 0001001011000000  
  715=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  716=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  717=>x"C043",	-- 1100000001000011  li	r3, 8
  718=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  719=>x"038B",	-- 0000001110001011  
  720=>x"D039",	-- 1101000000111001  lw	r1, r7
  721=>x"043F",	-- 0000010000111111  inc	r7, r7
  722=>x"D038",	-- 1101000000111000  lw	r0, r7
  723=>x"043F",	-- 0000010000111111  inc	r7, r7
  724=>x"0400",	-- 0000010000000000  inc	r0, r0
  725=>x"D03E",	-- 1101000000111110  lw	r6, r7
  726=>x"043F",	-- 0000010000111111  inc	r7, r7
  727=>x"E383",	-- 1110001110000011  ba	-, r6
  728=>x"063F",	-- 0000011000111111  dec	r7, r7
  729=>x"D23E",	-- 1101001000111110  sw	r6, r7
  730=>x"FFF4",	-- 1111111111110100  liw	r4, 10000
  731=>x"2710",	-- 0010011100010000  
  732=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  733=>x"02EB",	-- 0000001011101011  
  734=>x"FFF4",	-- 1111111111110100  liw	r4, 1000
  735=>x"03E8",	-- 0000001111101000  
  736=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  737=>x"02EB",	-- 0000001011101011  
  738=>x"C324",	-- 1100001100100100  li	r4, 100
  739=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  740=>x"02EB",	-- 0000001011101011  
  741=>x"C054",	-- 1100000001010100  li	r4, 10
  742=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  743=>x"02EB",	-- 0000001011101011  
  744=>x"D03E",	-- 1101000000111110  lw	r6, r7
  745=>x"043F",	-- 0000010000111111  inc	r7, r7
  746=>x"C00C",	-- 1100000000001100  li	r4, 1
  747=>x"C17B",	-- 1100000101111011  li	r3, 0x2F
  748=>x"041B",	-- 0000010000011011  inc	r3, r3
  749=>x"0B12",	-- 0000101100010010  sub	r2, r2, r4
  750=>x"BF91",	-- 1011111110010001  brige	r2, printnum.loop
  751=>x"0912",	-- 0000100100010010  add	r2, r2, r4
  752=>x"063F",	-- 0000011000111111  dec	r7, r7
  753=>x"D23E",	-- 1101001000111110  sw	r6, r7
  754=>x"063F",	-- 0000011000111111  dec	r7, r7
  755=>x"D23A",	-- 1101001000111010  sw	r2, r7
  756=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  757=>x"02C3",	-- 0000001011000011  
  758=>x"D03A",	-- 1101000000111010  lw	r2, r7
  759=>x"043F",	-- 0000010000111111  inc	r7, r7
  760=>x"D03E",	-- 1101000000111110  lw	r6, r7
  761=>x"043F",	-- 0000010000111111  inc	r7, r7
  762=>x"E383",	-- 1110001110000011  ba	-, r6
  763=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  764=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  765=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  766=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  767=>x"C0A0",	-- 1100000010100000  li	r0, 20
  768=>x"0412",	-- 0000010000010010  inc	r2, r2
  769=>x"D011",	-- 1101000000010001  lw	r1, r2
  770=>x"E421",	-- 1110010000100001  exw	r1, r4
  771=>x"0412",	-- 0000010000010010  inc	r2, r2
  772=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  773=>x"061B",	-- 0000011000011011  dec	r3, r3
  774=>x"BE9C",	-- 1011111010011100  brine	r3, put_sprite_16_aligned.loop
  775=>x"C005",	-- 1100000000000101  li	r5, 0
  776=>x"E383",	-- 1110001110000011  ba	-, r6
  777=>x"C07D",	-- 1100000001111101  li	r5, 15
  778=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  779=>x"6600",	-- 0110011000000000  shr	r0, r0, 3
  780=>x"BBE8",	-- 1011101111101000  brieq	r5, put_sprite_16_aligned
  781=>x"062D",	-- 0000011000101101  dec	r5, r5
  782=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  783=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  784=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  785=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  786=>x"063F",	-- 0000011000111111  dec	r7, r7
  787=>x"D23B",	-- 1101001000111011  sw	r3, r7
  788=>x"0412",	-- 0000010000010010  inc	r2, r2
  789=>x"D011",	-- 1101000000010001  lw	r1, r2
  790=>x"CFF8",	-- 1100111111111000  li	r0, -1
  791=>x"3D40",	-- 0011110101000000  rsr	r0, r0, r5
  792=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  793=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  794=>x"D023",	-- 1101000000100011  lw	r3, r4
  795=>x"2600",	-- 0010011000000000  not	r0, r0
  796=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  797=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  798=>x"E421",	-- 1110010000100001  exw	r1, r4
  799=>x"0424",	-- 0000010000100100  inc	r4, r4
  800=>x"D011",	-- 1101000000010001  lw	r1, r2
  801=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  802=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  803=>x"D023",	-- 1101000000100011  lw	r3, r4
  804=>x"2600",	-- 0010011000000000  not	r0, r0
  805=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  806=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  807=>x"E421",	-- 1110010000100001  exw	r1, r4
  808=>x"0412",	-- 0000010000010010  inc	r2, r2
  809=>x"C098",	-- 1100000010011000  li	r0, 19
  810=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  811=>x"D03B",	-- 1101000000111011  lw	r3, r7
  812=>x"043F",	-- 0000010000111111  inc	r7, r7
  813=>x"061B",	-- 0000011000011011  dec	r3, r3
  814=>x"B91C",	-- 1011100100011100  brine	r3, put_sprite_16.loop
  815=>x"C005",	-- 1100000000000101  li	r5, 0
  816=>x"E383",	-- 1110001110000011  ba	-, r6
  817=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  818=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  819=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  820=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  821=>x"C005",	-- 1100000000000101  li	r5, 0
  822=>x"D020",	-- 1101000000100000  lw	r0, r4
  823=>x"D011",	-- 1101000000010001  lw	r1, r2
  824=>x"0412",	-- 0000010000010010  inc	r2, r2
  825=>x"2040",	-- 0010000001000000  and	r0, r0, r1
  826=>x"D011",	-- 1101000000010001  lw	r1, r2
  827=>x"2240",	-- 0010001001000000  or	r0, r0, r1
  828=>x"E420",	-- 1110010000100000  exw	r0, r4
  829=>x"0612",	-- 0000011000010010  dec	r2, r2
  830=>x"D011",	-- 1101000000010001  lw	r1, r2
  831=>x"2609",	-- 0010011000001001  not	r1, r1
  832=>x"0412",	-- 0000010000010010  inc	r2, r2
  833=>x"2040",	-- 0010000001000000  and	r0, r0, r1
  834=>x"222D",	-- 0010001000101101  or	r5, r5, r0
  835=>x"0412",	-- 0000010000010010  inc	r2, r2
  836=>x"C0A0",	-- 1100000010100000  li	r0, 20
  837=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  838=>x"061B",	-- 0000011000011011  dec	r3, r3
  839=>x"AE5C",	-- 1010111001011100  brine	r3, put_sprite_16_aligned.loop
  840=>x"E383",	-- 1110001110000011  ba	-, r6
  841=>x"C07D",	-- 1100000001111101  li	r5, 15
  842=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  843=>x"6600",	-- 0110011000000000  shr	r0, r0, 3
  844=>x"B968",	-- 1011100101101000  brieq	r5, put_sprite_16_masked_aligned
  845=>x"062D",	-- 0000011000101101  dec	r5, r5
  846=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  847=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  848=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  849=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  850=>x"063F",	-- 0000011000111111  dec	r7, r7
  851=>x"D23E",	-- 1101001000111110  sw	r6, r7
  852=>x"102E",	-- 0001000000101110  mova	r6, r5
  853=>x"C005",	-- 1100000000000101  li	r5, 0
  854=>x"063F",	-- 0000011000111111  dec	r7, r7
  855=>x"D23B",	-- 1101001000111011  sw	r3, r7
  856=>x"063F",	-- 0000011000111111  dec	r7, r7
  857=>x"D23D",	-- 1101001000111101  sw	r5, r7
  858=>x"D010",	-- 1101000000010000  lw	r0, r2
  859=>x"3980",	-- 0011100110000000  rrr	r0, r0, r6
  860=>x"0412",	-- 0000010000010010  inc	r2, r2
  861=>x"D011",	-- 1101000000010001  lw	r1, r2
  862=>x"3989",	-- 0011100110001001  rrr	r1, r1, r6
  863=>x"CFFD",	-- 1100111111111101  li	r5, -1
  864=>x"3DAD",	-- 0011110110101101  rsr	r5, r5, r6
  865=>x"2149",	-- 0010000101001001  and	r1, r1, r5
  866=>x"D023",	-- 1101000000100011  lw	r3, r4
  867=>x"262D",	-- 0010011000101101  not	r5, r5
  868=>x"222D",	-- 0010001000101101  or	r5, r5, r0
  869=>x"215B",	-- 0010000101011011  and	r3, r3, r5
  870=>x"225B",	-- 0010001001011011  or	r3, r3, r1
  871=>x"E423",	-- 1110010000100011  exw	r3, r4
  872=>x"262D",	-- 0010011000101101  not	r5, r5
  873=>x"215B",	-- 0010000101011011  and	r3, r3, r5
  874=>x"D03D",	-- 1101000000111101  lw	r5, r7
  875=>x"043F",	-- 0000010000111111  inc	r7, r7
  876=>x"22ED",	-- 0010001011101101  or	r5, r5, r3
  877=>x"0424",	-- 0000010000100100  inc	r4, r4
  878=>x"063F",	-- 0000011000111111  dec	r7, r7
  879=>x"D23D",	-- 1101001000111101  sw	r5, r7
  880=>x"D011",	-- 1101000000010001  lw	r1, r2
  881=>x"3989",	-- 0011100110001001  rrr	r1, r1, r6
  882=>x"CFFD",	-- 1100111111111101  li	r5, -1
  883=>x"3DAD",	-- 0011110110101101  rsr	r5, r5, r6
  884=>x"262D",	-- 0010011000101101  not	r5, r5
  885=>x"2149",	-- 0010000101001001  and	r1, r1, r5
  886=>x"D023",	-- 1101000000100011  lw	r3, r4
  887=>x"262D",	-- 0010011000101101  not	r5, r5
  888=>x"222D",	-- 0010001000101101  or	r5, r5, r0
  889=>x"215B",	-- 0010000101011011  and	r3, r3, r5
  890=>x"225B",	-- 0010001001011011  or	r3, r3, r1
  891=>x"E423",	-- 1110010000100011  exw	r3, r4
  892=>x"262D",	-- 0010011000101101  not	r5, r5
  893=>x"215B",	-- 0010000101011011  and	r3, r3, r5
  894=>x"D03D",	-- 1101000000111101  lw	r5, r7
  895=>x"043F",	-- 0000010000111111  inc	r7, r7
  896=>x"22ED",	-- 0010001011101101  or	r5, r5, r3
  897=>x"0412",	-- 0000010000010010  inc	r2, r2
  898=>x"C098",	-- 1100000010011000  li	r0, 19
  899=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  900=>x"D03B",	-- 1101000000111011  lw	r3, r7
  901=>x"043F",	-- 0000010000111111  inc	r7, r7
  902=>x"061B",	-- 0000011000011011  dec	r3, r3
  903=>x"B3DC",	-- 1011001111011100  brine	r3, put_sprite_16_masked.loop
  904=>x"D03E",	-- 1101000000111110  lw	r6, r7
  905=>x"043F",	-- 0000010000111111  inc	r7, r7
  906=>x"E383",	-- 1110001110000011  ba	-, r6
  907=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  908=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  909=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  910=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  911=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  912=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  913=>x"C0A5",	-- 1100000010100101  li	r5, 20
  914=>x"8404",	-- 1000010000000100  brine	r0, put_sprite_8_aligned.loop1
  915=>x"D010",	-- 1101000000010000  lw	r0, r2
  916=>x"D021",	-- 1101000000100001  lw	r1, r4
  917=>x"1A41",	-- 0001101001000001  mixhl	r1, r0, r1
  918=>x"D221",	-- 1101001000100001  sw	r1, r4
  919=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  920=>x"061B",	-- 0000011000011011  dec	r3, r3
  921=>x"E398",	-- 1110001110011000  baeq	r3, r6
  922=>x"D021",	-- 1101000000100001  lw	r1, r4
  923=>x"1E41",	-- 0001111001000001  mixll	r1, r0, r1
  924=>x"D221",	-- 1101001000100001  sw	r1, r4
  925=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  926=>x"0412",	-- 0000010000010010  inc	r2, r2
  927=>x"061B",	-- 0000011000011011  dec	r3, r3
  928=>x"E398",	-- 1110001110011000  baeq	r3, r6
  929=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop0
  930=>x"D010",	-- 1101000000010000  lw	r0, r2
  931=>x"D021",	-- 1101000000100001  lw	r1, r4
  932=>x"1809",	-- 0001100000001001  mixhh	r1, r1, r0
  933=>x"D221",	-- 1101001000100001  sw	r1, r4
  934=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  935=>x"061B",	-- 0000011000011011  dec	r3, r3
  936=>x"E398",	-- 1110001110011000  baeq	r3, r6
  937=>x"D021",	-- 1101000000100001  lw	r1, r4
  938=>x"1A09",	-- 0001101000001001  mixhl	r1, r1, r0
  939=>x"D221",	-- 1101001000100001  sw	r1, r4
  940=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  941=>x"0412",	-- 0000010000010010  inc	r2, r2
  942=>x"061B",	-- 0000011000011011  dec	r3, r3
  943=>x"E398",	-- 1110001110011000  baeq	r3, r6
  944=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop1
  945=>x"C03D",	-- 1100000000111101  li	r5, 7
  946=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  947=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  948=>x"B5E8",	-- 1011010111101000  brieq	r5, put_sprite_8_aligned
  949=>x"062D",	-- 0000011000101101  dec	r5, r5
  950=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  951=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  952=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  953=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  954=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  955=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  956=>x"8A04",	-- 1000101000000100  brine	r0, put_sprite_8.loop1
  957=>x"D010",	-- 1101000000010000  lw	r0, r2
  958=>x"063F",	-- 0000011000111111  dec	r7, r7
  959=>x"D23A",	-- 1101001000111010  sw	r2, r7
  960=>x"C802",	-- 1100100000000010  li	r2, 0x100
  961=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  962=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  963=>x"D021",	-- 1101000000100001  lw	r1, r4
  964=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  965=>x"2612",	-- 0010011000010010  not	r2, r2
  966=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  967=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  968=>x"D221",	-- 1101001000100001  sw	r1, r4
  969=>x"C0A1",	-- 1100000010100001  li	r1, 20
  970=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  971=>x"D03A",	-- 1101000000111010  lw	r2, r7
  972=>x"043F",	-- 0000010000111111  inc	r7, r7
  973=>x"061B",	-- 0000011000011011  dec	r3, r3
  974=>x"E398",	-- 1110001110011000  baeq	r3, r6
  975=>x"D010",	-- 1101000000010000  lw	r0, r2
  976=>x"063F",	-- 0000011000111111  dec	r7, r7
  977=>x"D23A",	-- 1101001000111010  sw	r2, r7
  978=>x"1E00",	-- 0001111000000000  mixll	r0, r0, r0
  979=>x"C802",	-- 1100100000000010  li	r2, 0x100
  980=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  981=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  982=>x"D021",	-- 1101000000100001  lw	r1, r4
  983=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  984=>x"2612",	-- 0010011000010010  not	r2, r2
  985=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  986=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  987=>x"D221",	-- 1101001000100001  sw	r1, r4
  988=>x"C0A1",	-- 1100000010100001  li	r1, 20
  989=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  990=>x"D03A",	-- 1101000000111010  lw	r2, r7
  991=>x"043F",	-- 0000010000111111  inc	r7, r7
  992=>x"0412",	-- 0000010000010010  inc	r2, r2
  993=>x"061B",	-- 0000011000011011  dec	r3, r3
  994=>x"E398",	-- 1110001110011000  baeq	r3, r6
  995=>x"B683",	-- 1011011010000011  bri	-, put_sprite_8.loop0
  996=>x"D010",	-- 1101000000010000  lw	r0, r2
  997=>x"063F",	-- 0000011000111111  dec	r7, r7
  998=>x"D23A",	-- 1101001000111010  sw	r2, r7
  999=>x"063F",	-- 0000011000111111  dec	r7, r7
 1000=>x"D23B",	-- 1101001000111011  sw	r3, r7
 1001=>x"C802",	-- 1100100000000010  li	r2, 0x100
 1002=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
 1003=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
 1004=>x"2080",	-- 0010000010000000  and	r0, r0, r2
 1005=>x"D021",	-- 1101000000100001  lw	r1, r4
 1006=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
 1007=>x"261B",	-- 0010011000011011  not	r3, r3
 1008=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
 1009=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
 1010=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
 1011=>x"D221",	-- 1101001000100001  sw	r1, r4
 1012=>x"0424",	-- 0000010000100100  inc	r4, r4
 1013=>x"D021",	-- 1101000000100001  lw	r1, r4
 1014=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
 1015=>x"261B",	-- 0010011000011011  not	r3, r3
 1016=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
 1017=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
 1018=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
 1019=>x"D221",	-- 1101001000100001  sw	r1, r4
 1020=>x"C099",	-- 1100000010011001  li	r1, 19
 1021=>x"0864",	-- 0000100001100100  add	r4, r4, r1
 1022=>x"D03B",	-- 1101000000111011  lw	r3, r7
 1023=>x"043F",	-- 0000010000111111  inc	r7, r7
 1024=>x"D03A",	-- 1101000000111010  lw	r2, r7
 1025=>x"043F",	-- 0000010000111111  inc	r7, r7
 1026=>x"061B",	-- 0000011000011011  dec	r3, r3
 1027=>x"E398",	-- 1110001110011000  baeq	r3, r6
 1028=>x"D010",	-- 1101000000010000  lw	r0, r2
 1029=>x"4E00",	-- 0100111000000000  shl	r0, r0, 7
 1030=>x"063F",	-- 0000011000111111  dec	r7, r7
 1031=>x"D23A",	-- 1101001000111010  sw	r2, r7
 1032=>x"063F",	-- 0000011000111111  dec	r7, r7
 1033=>x"D23B",	-- 1101001000111011  sw	r3, r7
 1034=>x"C802",	-- 1100100000000010  li	r2, 0x100
 1035=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
 1036=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
 1037=>x"2080",	-- 0010000010000000  and	r0, r0, r2
 1038=>x"D021",	-- 1101000000100001  lw	r1, r4
 1039=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
 1040=>x"261B",	-- 0010011000011011  not	r3, r3
 1041=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
 1042=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
 1043=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
 1044=>x"D221",	-- 1101001000100001  sw	r1, r4
 1045=>x"0424",	-- 0000010000100100  inc	r4, r4
 1046=>x"D021",	-- 1101000000100001  lw	r1, r4
 1047=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
 1048=>x"261B",	-- 0010011000011011  not	r3, r3
 1049=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
 1050=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
 1051=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
 1052=>x"D221",	-- 1101001000100001  sw	r1, r4
 1053=>x"C099",	-- 1100000010011001  li	r1, 19
 1054=>x"0864",	-- 0000100001100100  add	r4, r4, r1
 1055=>x"D03B",	-- 1101000000111011  lw	r3, r7
 1056=>x"043F",	-- 0000010000111111  inc	r7, r7
 1057=>x"D03A",	-- 1101000000111010  lw	r2, r7
 1058=>x"043F",	-- 0000010000111111  inc	r7, r7
 1059=>x"0412",	-- 0000010000010010  inc	r2, r2
 1060=>x"061B",	-- 0000011000011011  dec	r3, r3
 1061=>x"E398",	-- 1110001110011000  baeq	r3, r6
 1062=>x"AF83",	-- 1010111110000011  bri	-, put_sprite_8.loop1
    others => x"0000"
    );
begin
  process(CLK)
  begin
    if (CLK'event AND CLK='1') then
      D <= m(to_integer(unsigned(AD)));
    end if;
  end process;
end Behavioral;
