----------------------------------------------------------------------------------
--
-- File retrieved, on 07/02/2010, from :
-- http://sebastien-viardot.imag.fr/Enseignements/Archi1A2s/sources/ROMPROG.vhd
--
-- Slightly altered to get rid of vendor-specific packages and adjust formatting
-- Now auto-filled by asrom script
--
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROMPROG is
  Port ( AD : in  STD_LOGIC_VECTOR (12 downto 0);
         D : out  STD_LOGIC_VECTOR (15 downto 0);
         CLK : in STD_LOGIC);
end ROMPROG;

architecture Behavioral of ROMPROG is
  constant low_address: natural := 0;
  constant high_address: natural := 8192;
  subtype octet is std_logic_vector( 15 downto 0 );
  type zone_memoire is
    array (natural range low_address to high_address-1) of octet;
  constant m: zone_memoire:= (
    0=>x"FFF7",	-- 1111111111110111  liw	r7, IRQ_mask
    1=>x"2000",	-- 0010000000000000  
    2=>x"F8C0",	-- 1111100011000000  bai	-, os_init
    3=>x"0100",	-- 0000000100000000  
   16=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_ack
   17=>x"2002",	-- 0010000000000010  
   18=>x"D001",	-- 1101000000000001  lw	r1, r0
   19=>x"F54A",	-- 1111010101001010  bspl	r2, r1, 5
   20=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_error
   21=>x"0050",	-- 0000000001010000  
   22=>x"F4CA",	-- 1111010011001010  bspl	r2, r1, 3
   23=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_kbd
   24=>x"0060",	-- 0000000001100000  
   25=>x"F40A",	-- 1111010000001010  bspl	r2, r1, 0
   26=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_tmr
   27=>x"0040",	-- 0000000001000000  
   28=>x"D201",	-- 1101001000000001  sw	r1, r0
   29=>x"FFFE",	-- 1111111111111110  reti
   64=>x"263F",	-- 0010011000111111  not r7, r7
   65=>x"D7C0",	-- 1101011111000000  out	r7
   66=>x"E383",	-- 1110001110000011  ba	-, r6
   80=>x"25FF",	-- 0010010111111111  xor	r7, r7, r7
   81=>x"D7C0",	-- 1101011111000000  out	r7
   82=>x"E383",	-- 1110001110000011  ba	-, r6
   96=>x"FFF2",	-- 1111111111110010  liw	r2, PS2_rx
   97=>x"2004",	-- 0010000000000100  
   98=>x"D012",	-- 1101000000010010  lw	r2, r2
   99=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map + 8
  100=>x"16C8",	-- 0001011011001000  
  101=>x"D01B",	-- 1101000000011011  lw	r3, r3
  102=>x"1EBF",	-- 0001111010111111  mixll	r7, r7, r2
  103=>x"C784",	-- 1100011110000100  li	r4, 0xF0
  104=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  105=>x"8B20",	-- 1000101100100000  brieq	r4, int_kbd.release
  106=>x"C704",	-- 1100011100000100  li	r4, 0xE0
  107=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  108=>x"88E0",	-- 1000100011100000  brieq	r4, int_kbd.extended
  109=>x"FFF5",	-- 1111111111110101  liw	r5, paper_keys - 1
  110=>x"16CF",	-- 0001011011001111  
  111=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  112=>x"80E0",	-- 1000000011100000  brieq	r4, $+3
  113=>x"FFF5",	-- 1111111111110101  liw	r5, paper_keys + 11 - 1
  114=>x"16DA",	-- 0001011011011010  
  115=>x"042D",	-- 0000010000101101  inc	r5, r5
  116=>x"D02C",	-- 1101000000101100  lw	r4, r5
  117=>x"8560",	-- 1000010101100000  brieq	r4, scan_code_mismatch
  118=>x"6E24",	-- 0110111000100100  shr	r4, r4, 7
  119=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  120=>x"BEE4",	-- 1011111011100100  brine	r4, scan_code_loop
  121=>x"D02A",	-- 1101000000101010  lw	r2, r5
  122=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  123=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  124=>x"741B",	-- 0111010000011011  shr	r3, r3, 10
  125=>x"C00D",	-- 1100000000001101  li	r5, 1
  126=>x"0612",	-- 0000011000010010  dec	r2, r2
  127=>x"3AAA",	-- 0011101010101010  rrl	r2, r5, r2
  128=>x"FFF5",	-- 1111111111110101  liw	r5, key_press_map
  129=>x"16C0",	-- 0001011011000000  
  130=>x"08ED",	-- 0000100011101101  add	r5, r5, r3
  131=>x"D02B",	-- 1101000000101011  lw	r3, r5
  132=>x"80E4",	-- 1000000011100100  brine	r4, scan_code_release
  133=>x"229B",	-- 0010001010011011  or	r3, r3, r2
  134=>x"80C3",	-- 1000000011000011  bri	-, scan_code_notify
  135=>x"2612",	-- 0010011000010010  not	r2, r2
  136=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  137=>x"D22B",	-- 1101001000101011  sw	r3, r5
  138=>x"C003",	-- 1100000000000011  li	r3, 0
  139=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  140=>x"16C8",	-- 0001011011001000  
  141=>x"D223",	-- 1101001000100011  sw	r3, r4
  142=>x"E383",	-- 1110001110000011  ba	-, r6
  143=>x"C014",	-- 1100000000010100  li	r4, 2
  144=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  145=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  146=>x"16C8",	-- 0001011011001000  
  147=>x"D223",	-- 1101001000100011  sw	r3, r4
  148=>x"E383",	-- 1110001110000011  ba	-, r6
  149=>x"C00C",	-- 1100000000001100  li	r4, 1
  150=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  151=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  152=>x"16C8",	-- 0001011011001000  
  153=>x"D223",	-- 1101001000100011  sw	r3, r4
  154=>x"E383",	-- 1110001110000011  ba	-, r6
  256=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_mask
  257=>x"2000",	-- 0010000000000000  
  258=>x"C0C9",	-- 1100000011001001  li	r1, 0x19
  259=>x"D201",	-- 1101001000000001  sw	r1, r0
  260=>x"0400",	-- 0000010000000000  inc	r0, r0
  261=>x"CFF9",	-- 1100111111111001  li	r1, -1
  262=>x"D201",	-- 1101001000000001  sw	r1, r0
  263=>x"C03A",	-- 1100000000111010  li	r2, 7
  264=>x"0880",	-- 0000100010000000  add	r0, r0, r2
  265=>x"C0EA",	-- 1100000011101010  li	r2, 0x1D
  266=>x"D202",	-- 1101001000000010  sw	r2, r0
  267=>x"0400",	-- 0000010000000000  inc	r0, r0
  268=>x"C07A",	-- 1100000001111010  li	r2, 15
  269=>x"D202",	-- 1101001000000010  sw	r2, r0
  270=>x"0400",	-- 0000010000000000  inc	r0, r0
  271=>x"C0DA",	-- 1100000011011010  li	r2, 0x1B
  272=>x"D202",	-- 1101001000000010  sw	r2, r0
  273=>x"0400",	-- 0000010000000000  inc	r0, r0
  274=>x"FFF2",	-- 1111111111110010  liw	r2, 817
  275=>x"0331",	-- 0000001100110001  
  276=>x"D202",	-- 1101001000000010  sw	r2, r0
  277=>x"FFF0",	-- 1111111111110000  liw	r0, key_press_map
  278=>x"16C0",	-- 0001011011000000  
  279=>x"C001",	-- 1100000000000001  li	r1, 0
  280=>x"C042",	-- 1100000001000010  li	r2, 8
  281=>x"D201",	-- 1101001000000001  sw	r1, r0
  282=>x"0400",	-- 0000010000000000  inc	r0, r0
  283=>x"0612",	-- 0000011000010010  dec	r2, r2
  284=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  285=>x"C0F3",	-- 1100000011110011  li	r3, 30
  286=>x"CFFA",	-- 1100111111111010  li	r2, -1
  287=>x"D21A",	-- 1101001000011010  sw	r2, r3
  288=>x"8083",	-- 1000000010000011  bri	-, PaperGameStart
  289=>x"8003",	-- 1000000000000011  bri	-, PaperMenuLoop
  290=>x"FFF0",	-- 1111111111110000  liw	r0, paper_dir
  291=>x"179C",	-- 0001011110011100  
  292=>x"C001",	-- 1100000000000001  li	r1, 0
  293=>x"D201",	-- 1101001000000001  sw	r1, r0
  294=>x"0400",	-- 0000010000000000  inc	r0, r0
  295=>x"FFF1",	-- 1111111111110001  liw	r1, 152 * 8
  296=>x"04C0",	-- 0000010011000000  
  297=>x"D201",	-- 1101001000000001  sw	r1, r0
  298=>x"0400",	-- 0000010000000000  inc	r0, r0
  299=>x"C001",	-- 1100000000000001  li	r1, 0
  300=>x"D201",	-- 1101001000000001  sw	r1, r0
  301=>x"0400",	-- 0000010000000000  inc	r0, r0
  302=>x"FFF1",	-- 1111111111110001  liw	r1, 128 * 8
  303=>x"0400",	-- 0000010000000000  
  304=>x"D201",	-- 1101001000000001  sw	r1, r0
  305=>x"0400",	-- 0000010000000000  inc	r0, r0
  306=>x"C001",	-- 1100000000000001  li	r1, 0
  307=>x"D201",	-- 1101001000000001  sw	r1, r0
  308=>x"0400",	-- 0000010000000000  inc	r0, r0
  309=>x"C069",	-- 1100000001101001  li	r1, 13
  310=>x"D201",	-- 1101001000000001  sw	r1, r0
  311=>x"0400",	-- 0000010000000000  inc	r0, r0
  312=>x"C011",	-- 1100000000010001  li	r1, 2
  313=>x"D201",	-- 1101001000000001  sw	r1, r0
  314=>x"0400",	-- 0000010000000000  inc	r0, r0
  315=>x"CFF8",	-- 1100111111111000  li	r0, -1
  316=>x"FAC6",	-- 1111101011000110  bail	-, r6, rand16_init
  317=>x"0243",	-- 0000001001000011  
  318=>x"C000",	-- 1100000000000000  li	r0, 0
  319=>x"CFF9",	-- 1100111111111001  li	r1, -1
  320=>x"C0A2",	-- 1100000010100010  li	r2, 20
  321=>x"D201",	-- 1101001000000001  sw	r1, r0
  322=>x"0400",	-- 0000010000000000  inc	r0, r0
  323=>x"0612",	-- 0000011000010010  dec	r2, r2
  324=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  325=>x"C001",	-- 1100000000000001  li	r1, 0
  326=>x"FFF2",	-- 1111111111110010  liw	r2, 18*20
  327=>x"0168",	-- 0000000101101000  
  328=>x"D201",	-- 1101001000000001  sw	r1, r0
  329=>x"0400",	-- 0000010000000000  inc	r0, r0
  330=>x"0612",	-- 0000011000010010  dec	r2, r2
  331=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  332=>x"CFF9",	-- 1100111111111001  li	r1, -1
  333=>x"C0A2",	-- 1100000010100010  li	r2, 20
  334=>x"D201",	-- 1101001000000001  sw	r1, r0
  335=>x"0400",	-- 0000010000000000  inc	r0, r0
  336=>x"0612",	-- 0000011000010010  dec	r2, r2
  337=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  338=>x"C020",	-- 1100000000100000  li	r0, 4
  339=>x"C029",	-- 1100000000101001  li	r1, 5
  340=>x"FFF2",	-- 1111111111110010  liw	r2, paper_title
  341=>x"17A4",	-- 0001011110100100  
  342=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  343=>x"0289",	-- 0000001010001001  
  344=>x"C778",	-- 1100011101111000  li	r0, 239
  345=>x"C009",	-- 1100000000001001  li	r1, 1
  346=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud
  347=>x"1780",	-- 0001011110000000  
  348=>x"C043",	-- 1100000001000011  li	r3, 8
  349=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  350=>x"0391",	-- 0000001110010001  
  351=>x"C0F8",	-- 1100000011111000  li	r0, 31
  352=>x"C009",	-- 1100000000001001  li	r1, 1
  353=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed + 1
  354=>x"17A1",	-- 0001011110100001  
  355=>x"D012",	-- 1101000000010010  lw	r2, r2
  356=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum
  357=>x"02B8",	-- 0000001010111000  
  358=>x"C120",	-- 1100000100100000  li	r0, 36
  359=>x"C009",	-- 1100000000001001  li	r1, 1
  360=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  361=>x"17AA",	-- 0001011110101010  
  362=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  363=>x"0289",	-- 0000001010001001  
  364=>x"C778",	-- 1100011101111000  li	r0, 239
  365=>x"C051",	-- 1100000001010001  li	r1, 10
  366=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud + 4
  367=>x"1784",	-- 0001011110000100  
  368=>x"C043",	-- 1100000001000011  li	r3, 8
  369=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  370=>x"0391",	-- 0000001110010001  
  371=>x"C0F8",	-- 1100000011111000  li	r0, 31
  372=>x"C051",	-- 1100000001010001  li	r1, 10
  373=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed + 2
  374=>x"17A2",	-- 0001011110100010  
  375=>x"D012",	-- 1101000000010010  lw	r2, r2
  376=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum
  377=>x"02B8",	-- 0000001010111000  
  378=>x"C120",	-- 1100000100100000  li	r0, 36
  379=>x"C051",	-- 1100000001010001  li	r1, 10
  380=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  381=>x"17AA",	-- 0001011110101010  
  382=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  383=>x"0289",	-- 0000001010001001  
  384=>x"FFF0",	-- 1111111111110000  liw	r0, 20*20
  385=>x"0190",	-- 0000000110010000  
  386=>x"C001",	-- 1100000000000001  li	r1, 0
  387=>x"FFF2",	-- 1111111111110010  liw	r2, 220*20
  388=>x"1130",	-- 0001000100110000  
  389=>x"D201",	-- 1101001000000001  sw	r1, r0
  390=>x"0400",	-- 0000010000000000  inc	r0, r0
  391=>x"0612",	-- 0000011000010010  dec	r2, r2
  392=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  393=>x"FFF5",	-- 1111111111110101  liw	r5, paper_tilemap
  394=>x"17B0",	-- 0001011110110000  
  395=>x"D02C",	-- 1101000000101100  lw	r4, r5
  396=>x"042D",	-- 0000010000101101  inc	r5, r5
  397=>x"8960",	-- 1000100101100000  brieq	r4, PaperGameTileSkip
  398=>x"063F",	-- 0000011000111111  dec	r7, r7
  399=>x"D23D",	-- 1101001000111101  sw	r5, r7
  400=>x"FFF3",	-- 1111111111110011  liw	r3, paper_tilemap
  401=>x"17B0",	-- 0001011110110000  
  402=>x"0AEB",	-- 0000101011101011  sub	r3, r5, r3
  403=>x"6E20",	-- 0110111000100000  shr	r0, r4, 7
  404=>x"6219",	-- 0110001000011001  shr	r1, r3, 1
  405=>x"4809",	-- 0100100000001001  shl	r1, r1, 4
  406=>x"C19A",	-- 1100000110011010  li	r2, 51
  407=>x"0889",	-- 0000100010001001  add	r1, r1, r2
  408=>x"FFF2",	-- 1111111111110010  liw	r2, paper_pos + 1
  409=>x"179E",	-- 0001011110011110  
  410=>x"D012",	-- 1101000000010010  lw	r2, r2
  411=>x"6412",	-- 0110010000010010  shr	r2, r2, 2
  412=>x"C0FB",	-- 1100000011111011  li	r3, 31
  413=>x"20D2",	-- 0010000011010010  and	r2, r2, r3
  414=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  415=>x"4E24",	-- 0100111000100100  shl	r4, r4, 7
  416=>x"6E24",	-- 0110111000100100  shr	r4, r4, 7
  417=>x"C00B",	-- 1100000000001011  li	r3, 1
  418=>x"FB06",	-- 1111101100000110  bailne	r0, r6, put_tile
  419=>x"0259",	-- 0000001001011001  
  420=>x"81E0",	-- 1000000111100000  brieq	r4, PaperGameSegmentSkip
  422=>x"C013",	-- 1100000000010011  li	r3, 2
  423=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_tile
  424=>x"0259",	-- 0000001001011001  
  425=>x"0624",	-- 0000011000100100  dec	r4, r4
  426=>x"BF64",	-- 1011111101100100  brine	r4, PaperGameSegmentLoop
  427=>x"C003",	-- 1100000000000011  li	r3, 0
  428=>x"C144",	-- 1100000101000100  li	r4, 40
  429=>x"0B04",	-- 0000101100000100  sub	r4, r0, r4
  430=>x"FB66",	-- 1111101101100110  baillt	r4, r6, put_tile
  431=>x"0259",	-- 0000001001011001  
  432=>x"D03D",	-- 1101000000111101  lw	r5, r7
  433=>x"043F",	-- 0000010000111111  inc	r7, r7
  434=>x"FFF4",	-- 1111111111110100  liw r4, paper_tilemap + 24
  435=>x"17C8",	-- 0001011111001000  
  436=>x"0B2C",	-- 0000101100101100  sub	r4, r5, r4
  437=>x"B5A5",	-- 1011010110100101  brilt	r4, PaperGameTileLoop
  438=>x"FFF3",	-- 1111111111110011  liw	r3, paper_speed
  439=>x"17A0",	-- 0001011110100000  
  440=>x"D01B",	-- 1101000000011011  lw	r3, r3
  441=>x"CFC4",	-- 1100111111000100  li	r4, 0x1F8
  442=>x"211C",	-- 0010000100011100  and	r4, r3, r4
  443=>x"0924",	-- 0000100100100100  add	r4, r4, r4
  444=>x"0924",	-- 0000100100100100  add	r4, r4, r4
  445=>x"FFF3",	-- 1111111111110011  liw	r3, paper_pos
  446=>x"179D",	-- 0001011110011101  
  447=>x"D018",	-- 1101000000011000  lw	r0, r3
  448=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  449=>x"FFF2",	-- 1111111111110010  liw	r2, paper_sprites
  450=>x"1720",	-- 0001011100100000  
  451=>x"0912",	-- 0000100100010010  add	r2, r2, r4
  452=>x"C161",	-- 1100000101100001  li	r1, 44
  453=>x"C083",	-- 1100000010000011  li	r3, 16
  454=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_16_masked
  455=>x"0329",	-- 0000001100101001  
  456=>x"906C",	-- 1001000001101100  brine	r5, PaperGameFail
  458=>x"C028",	-- 1100000000101000  li	r0, 5
  459=>x"C001",	-- 1100000000000001  li	r1, 0
  460=>x"8043",	-- 1000000001000011  bri	-, $+1
  461=>x"0609",	-- 0000011000001001  dec	r1, r1
  462=>x"BF8C",	-- 1011111110001100  brine	r1, $-2
  463=>x"0600",	-- 0000011000000000  dec	r0, r0
  464=>x"BEC4",	-- 1011111011000100  brine	r0, $-5
  465=>x"FFF2",	-- 1111111111110010  liw	r2, paper_pos
  466=>x"179D",	-- 0001011110011101  
  467=>x"FFF3",	-- 1111111111110011  liw	r3, paper_speed
  468=>x"17A0",	-- 0001011110100000  
  469=>x"D010",	-- 1101000000010000  lw	r0, r2
  470=>x"D019",	-- 1101000000011001  lw	r1, r3
  471=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  472=>x"8C45",	-- 1000110001000101  brilt	r0, PaperGameFail
  473=>x"FFF4",	-- 1111111111110100  liw	r4, 304*8
  474=>x"0980",	-- 0000100110000000  
  475=>x"0B04",	-- 0000101100000100  sub	r4, r0, r4
  476=>x"8B61",	-- 1000101101100001  brige	r4, PaperGameFail
  477=>x"D210",	-- 1101001000010000  sw	r0, r2
  478=>x"0412",	-- 0000010000010010  inc	r2, r2
  479=>x"041B",	-- 0000010000011011  inc	r3, r3
  480=>x"D010",	-- 1101000000010000  lw	r0, r2
  481=>x"D019",	-- 1101000000011001  lw	r1, r3
  482=>x"C7FC",	-- 1100011111111100  li	r4, 0xFF
  483=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  484=>x"2101",	-- 0010000100000001  and	r1, r0, r4
  485=>x"D211",	-- 1101001000010001  sw	r1, r2
  486=>x"2624",	-- 0010011000100100  not	r4, r4
  487=>x"2100",	-- 0010000100000000  and	r0, r0, r4
  488=>x"FB06",	-- 1111101100000110  bailne	r0, r6, PaperMapScroll
  489=>x"0217",	-- 0000001000010111  
  490=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  491=>x"16C0",	-- 0001011011000000  
  492=>x"D01B",	-- 1101000000011011  lw	r3, r3
  493=>x"F818",	-- 1111100000011000  baieq	r3, PaperGameRedrawContent
  494=>x"0180",	-- 0000000110000000  
  495=>x"F7DC",	-- 1111011111011100  bspl	r4, r3, 15
  496=>x"89A4",	-- 1000100110100100  brine	r4, PaperGameQuit
  497=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  498=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveUp
  499=>x"F49C",	-- 1111010010011100  bspl	r4, r3, 2
  500=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveDOWN
  501=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  502=>x"8220",	-- 1000001000100000  brieq	r4, PaperNoMoveLEFT
  503=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  504=>x"17A0",	-- 0001011110100000  
  505=>x"D010",	-- 1101000000010000  lw	r0, r2
  506=>x"0600",	-- 0000011000000000  dec	r0, r0
  507=>x"0600",	-- 0000011000000000  dec	r0, r0
  508=>x"0600",	-- 0000011000000000  dec	r0, r0
  509=>x"D210",	-- 1101001000010000  sw	r0, r2
  510=>x"F4DC",	-- 1111010011011100  bspl	r4, r3, 3
  511=>x"8220",	-- 1000001000100000  brieq	r4, PaperNoMoveRIGHT
  512=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  513=>x"17A0",	-- 0001011110100000  
  514=>x"D010",	-- 1101000000010000  lw	r0, r2
  515=>x"0400",	-- 0000010000000000  inc	r0, r0
  516=>x"0400",	-- 0000010000000000  inc	r0, r0
  517=>x"0400",	-- 0000010000000000  inc	r0, r0
  518=>x"D210",	-- 1101001000010000  sw	r0, r2
  519=>x"F8C0",	-- 1111100011000000  bai	-, PaperGameRedrawContent
  520=>x"0180",	-- 0000000110000000  
  521=>x"C000",	-- 1100000000000000  li	r0, 0
  522=>x"FFF2",	-- 1111111111110010  liw	r2, 240*20
  523=>x"12C0",	-- 0001001011000000  
  524=>x"D001",	-- 1101000000000001  lw	r1, r0
  525=>x"2609",	-- 0010011000001001  not	r1, r1
  526=>x"D201",	-- 1101001000000001  sw	r1, r0
  527=>x"0400",	-- 0000010000000000  inc	r0, r0
  528=>x"0612",	-- 0000011000010010  dec	r2, r2
  529=>x"BED4",	-- 1011111011010100  brine	r2, $-5
  530=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  531=>x"16C0",	-- 0001011011000000  
  532=>x"D01A",	-- 1101000000011010  lw	r2, r3
  533=>x"BFD0",	-- 1011111111010000  brieq	r2, $-1
  534=>x"FFFF",	-- 1111111111111111  reset
  535=>x"FFF0",	-- 1111111111110000  liw	r0, paper_tilemap
  536=>x"17B0",	-- 0001011110110000  
  537=>x"C021",	-- 1100000000100001  li	r1, 4
  538=>x"0841",	-- 0000100001000001  add	r1, r0, r1
  539=>x"C0A2",	-- 1100000010100010  li	r2, 5*4
  540=>x"D00B",	-- 1101000000001011  lw	r3, r1
  541=>x"D203",	-- 1101001000000011  sw	r3, r0
  542=>x"0400",	-- 0000010000000000  inc	r0, r0
  543=>x"0409",	-- 0000010000001001  inc	r1, r1
  544=>x"0612",	-- 0000011000010010  dec	r2, r2
  545=>x"BED4",	-- 1011111011010100  brine	r2, PaperGameScrollLoop
  546=>x"063F",	-- 0000011000111111  dec	r7, r7
  547=>x"D23E",	-- 1101001000111110  sw	r6, r7
  548=>x"FAC6",	-- 1111101011000110  bail	-, r6, rand16
  549=>x"0247",	-- 0000001001000111  
  550=>x"C03A",	-- 1100000000111010  li	r2, 0x07
  551=>x"208B",	-- 0010000010001011  and	r3, r1, r2
  552=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  553=>x"208C",	-- 0010000010001100  and	r4, r1, r2
  554=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  555=>x"1F19",	-- 0001111100011001  mixll	r1, r3, r4
  556=>x"D201",	-- 1101001000000001  sw	r1, r0
  557=>x"0400",	-- 0000010000000000  inc	r0, r0
  558=>x"091C",	-- 0000100100011100  add r4, r3, r4
  559=>x"208B",	-- 0010000010001011  and	r3, r1, r2
  560=>x"091C",	-- 0000100100011100  add r4, r3, r4
  561=>x"0424",	-- 0000010000100100  inc	r4, r4
  562=>x"6209",	-- 0110001000001001  shr	r1, r1, 1
  563=>x"208B",	-- 0010000010001011  and	r3, r1, r2
  564=>x"091B",	-- 0000100100011011  add r3, r3, r4
  565=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  566=>x"208C",	-- 0010000010001100  and	r4, r1, r2
  567=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  568=>x"1F19",	-- 0001111100011001  mixll	r1, r3, r4
  569=>x"D201",	-- 1101001000000001  sw	r1, r0
  570=>x"0400",	-- 0000010000000000  inc	r0, r0
  571=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed + 1
  572=>x"17A1",	-- 0001011110100001  
  573=>x"D011",	-- 1101000000010001  lw	r1, r2
  574=>x"0409",	-- 0000010000001001  inc	r1, r1
  575=>x"D211",	-- 1101001000010001  sw	r1, r2
  576=>x"D03E",	-- 1101000000111110  lw	r6, r7
  577=>x"043F",	-- 0000010000111111  inc	r7, r7
  578=>x"E383",	-- 1110001110000011  ba	-, r6
  579=>x"FFF2",	-- 1111111111110010  liw	r2, rand_seed
  580=>x"16C8",	-- 0001011011001000  
  581=>x"D210",	-- 1101001000010000  sw	r0, r2
  582=>x"E383",	-- 1110001110000011  ba	-, r6
  583=>x"FFF2",	-- 1111111111110010  liw	r2, rand_seed
  584=>x"16C8",	-- 0001011011001000  
  585=>x"D013",	-- 1101000000010011  lw	r3, r2
  586=>x"C7EC",	-- 1100011111101100  li	r4, 253
  587=>x"1F19",	-- 0001111100011001  mixll	r1, r3, r4
  588=>x"18E4",	-- 0001100011100100  mixhh	r4, r4, r3
  589=>x"C002",	-- 1100000000000010  li	r2, 0
  590=>x"0AC9",	-- 0000101011001001  sub	r1, r1, r3
  591=>x"0EA4",	-- 0000111010100100  sbc	r4, r4, r2
  592=>x"0EC9",	-- 0000111011001001  sbc	r1, r1, r3
  593=>x"0EA4",	-- 0000111010100100  sbc	r4, r4, r2
  594=>x"1B13",	-- 0001101100010011  mixhl	r3, r2, r4
  595=>x"0EC9",	-- 0000111011001001  sbc	r1, r1, r3
  596=>x"0C89",	-- 0000110010001001  adc	r1, r1, r2
  597=>x"FFF2",	-- 1111111111110010  liw	r2, rand_seed
  598=>x"16C8",	-- 0001011011001000  
  599=>x"D211",	-- 1101001000010001  sw	r1, r2
  600=>x"E383",	-- 1110001110000011  ba	-, r6
  601=>x"063F",	-- 0000011000111111  dec	r7, r7
  602=>x"D238",	-- 1101001000111000  sw	r0, r7
  603=>x"063F",	-- 0000011000111111  dec	r7, r7
  604=>x"D239",	-- 1101001000111001  sw	r1, r7
  605=>x"063F",	-- 0000011000111111  dec	r7, r7
  606=>x"D23A",	-- 1101001000111010  sw	r2, r7
  607=>x"063F",	-- 0000011000111111  dec	r7, r7
  608=>x"D23B",	-- 1101001000111011  sw	r3, r7
  609=>x"063F",	-- 0000011000111111  dec	r7, r7
  610=>x"D23C",	-- 1101001000111100  sw	r4, r7
  611=>x"063F",	-- 0000011000111111  dec	r7, r7
  612=>x"D23D",	-- 1101001000111101  sw	r5, r7
  613=>x"063F",	-- 0000011000111111  dec	r7, r7
  614=>x"D23E",	-- 1101001000111110  sw	r6, r7
  615=>x"FFF2",	-- 1111111111110010  liw	r2, paper_tiles
  616=>x"1790",	-- 0001011110010000  
  617=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  618=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  619=>x"C043",	-- 1100000001000011  li	r3, 8
  620=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  621=>x"036B",	-- 0000001101101011  
  622=>x"D03E",	-- 1101000000111110  lw	r6, r7
  623=>x"043F",	-- 0000010000111111  inc	r7, r7
  624=>x"D03D",	-- 1101000000111101  lw	r5, r7
  625=>x"043F",	-- 0000010000111111  inc	r7, r7
  626=>x"D03C",	-- 1101000000111100  lw	r4, r7
  627=>x"043F",	-- 0000010000111111  inc	r7, r7
  628=>x"D03B",	-- 1101000000111011  lw	r3, r7
  629=>x"043F",	-- 0000010000111111  inc	r7, r7
  630=>x"D03A",	-- 1101000000111010  lw	r2, r7
  631=>x"043F",	-- 0000010000111111  inc	r7, r7
  632=>x"D039",	-- 1101000000111001  lw	r1, r7
  633=>x"043F",	-- 0000010000111111  inc	r7, r7
  634=>x"D038",	-- 1101000000111000  lw	r0, r7
  635=>x"043F",	-- 0000010000111111  inc	r7, r7
  636=>x"0400",	-- 0000010000000000  inc	r0, r0
  637=>x"E383",	-- 1110001110000011  ba	-, r6
  638=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  639=>x"C084",	-- 1100000010000100  li	r4, 16
  640=>x"0800",	-- 0000100000000000  add	r0, r0, r0
  641=>x"0C49",	-- 0000110001001001  adc	r1, r1, r1
  642=>x"0A8B",	-- 0000101010001011  sub	r3, r1, r2
  643=>x"80DD",	-- 1000000011011101  brilt	r3, div_16_16.skip
  644=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  645=>x"0400",	-- 0000010000000000  inc	r0, r0
  646=>x"0624",	-- 0000011000100100  dec	r4, r4
  647=>x"BE64",	-- 1011111001100100  brine	r4, div_16_16.loop
  648=>x"E383",	-- 1110001110000011  ba	-, r6
  649=>x"063F",	-- 0000011000111111  dec	r7, r7
  650=>x"D23E",	-- 1101001000111110  sw	r6, r7
  651=>x"D013",	-- 1101000000010011  lw	r3, r2
  652=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  653=>x"84D8",	-- 1000010011011000  brieq	r3, puts.end
  654=>x"063F",	-- 0000011000111111  dec	r7, r7
  655=>x"D23A",	-- 1101001000111010  sw	r2, r7
  656=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  657=>x"02A3",	-- 0000001010100011  
  658=>x"D03A",	-- 1101000000111010  lw	r2, r7
  659=>x"043F",	-- 0000010000111111  inc	r7, r7
  660=>x"D013",	-- 1101000000010011  lw	r3, r2
  661=>x"4E1B",	-- 0100111000011011  shl	r3, r3, 7
  662=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  663=>x"8258",	-- 1000001001011000  brieq	r3, puts.end
  664=>x"063F",	-- 0000011000111111  dec	r7, r7
  665=>x"D23A",	-- 1101001000111010  sw	r2, r7
  666=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  667=>x"02A3",	-- 0000001010100011  
  668=>x"D03A",	-- 1101000000111010  lw	r2, r7
  669=>x"043F",	-- 0000010000111111  inc	r7, r7
  670=>x"0412",	-- 0000010000010010  inc	r2, r2
  671=>x"BB03",	-- 1011101100000011  bri	-, puts.loop
  672=>x"D03E",	-- 1101000000111110  lw	r6, r7
  673=>x"043F",	-- 0000010000111111  inc	r7, r7
  674=>x"E383",	-- 1110001110000011  ba	-, r6
  675=>x"063F",	-- 0000011000111111  dec	r7, r7
  676=>x"D23E",	-- 1101001000111110  sw	r6, r7
  677=>x"063F",	-- 0000011000111111  dec	r7, r7
  678=>x"D238",	-- 1101001000111000  sw	r0, r7
  679=>x"063F",	-- 0000011000111111  dec	r7, r7
  680=>x"D239",	-- 1101001000111001  sw	r1, r7
  681=>x"FFF2",	-- 1111111111110010  liw	r2, font_map
  682=>x"12C0",	-- 0001001011000000  
  683=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  684=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  685=>x"C043",	-- 1100000001000011  li	r3, 8
  686=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  687=>x"036B",	-- 0000001101101011  
  688=>x"D039",	-- 1101000000111001  lw	r1, r7
  689=>x"043F",	-- 0000010000111111  inc	r7, r7
  690=>x"D038",	-- 1101000000111000  lw	r0, r7
  691=>x"043F",	-- 0000010000111111  inc	r7, r7
  692=>x"0400",	-- 0000010000000000  inc	r0, r0
  693=>x"D03E",	-- 1101000000111110  lw	r6, r7
  694=>x"043F",	-- 0000010000111111  inc	r7, r7
  695=>x"E383",	-- 1110001110000011  ba	-, r6
  696=>x"063F",	-- 0000011000111111  dec	r7, r7
  697=>x"D23E",	-- 1101001000111110  sw	r6, r7
  698=>x"FFF4",	-- 1111111111110100  liw	r4, 10000
  699=>x"2710",	-- 0010011100010000  
  700=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  701=>x"02CB",	-- 0000001011001011  
  702=>x"FFF4",	-- 1111111111110100  liw	r4, 1000
  703=>x"03E8",	-- 0000001111101000  
  704=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  705=>x"02CB",	-- 0000001011001011  
  706=>x"C324",	-- 1100001100100100  li	r4, 100
  707=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  708=>x"02CB",	-- 0000001011001011  
  709=>x"C054",	-- 1100000001010100  li	r4, 10
  710=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  711=>x"02CB",	-- 0000001011001011  
  712=>x"D03E",	-- 1101000000111110  lw	r6, r7
  713=>x"043F",	-- 0000010000111111  inc	r7, r7
  714=>x"C00C",	-- 1100000000001100  li	r4, 1
  715=>x"C17B",	-- 1100000101111011  li	r3, 0x2F
  716=>x"041B",	-- 0000010000011011  inc	r3, r3
  717=>x"0B12",	-- 0000101100010010  sub	r2, r2, r4
  718=>x"BF91",	-- 1011111110010001  brige	r2, printnum.loop
  719=>x"0912",	-- 0000100100010010  add	r2, r2, r4
  720=>x"063F",	-- 0000011000111111  dec	r7, r7
  721=>x"D23E",	-- 1101001000111110  sw	r6, r7
  722=>x"063F",	-- 0000011000111111  dec	r7, r7
  723=>x"D23A",	-- 1101001000111010  sw	r2, r7
  724=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  725=>x"02A3",	-- 0000001010100011  
  726=>x"D03A",	-- 1101000000111010  lw	r2, r7
  727=>x"043F",	-- 0000010000111111  inc	r7, r7
  728=>x"D03E",	-- 1101000000111110  lw	r6, r7
  729=>x"043F",	-- 0000010000111111  inc	r7, r7
  730=>x"E383",	-- 1110001110000011  ba	-, r6
  731=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  732=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  733=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  734=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  735=>x"C0A0",	-- 1100000010100000  li	r0, 20
  736=>x"0412",	-- 0000010000010010  inc	r2, r2
  737=>x"D011",	-- 1101000000010001  lw	r1, r2
  738=>x"E421",	-- 1110010000100001  exw	r1, r4
  739=>x"0412",	-- 0000010000010010  inc	r2, r2
  740=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  741=>x"061B",	-- 0000011000011011  dec	r3, r3
  742=>x"BE9C",	-- 1011111010011100  brine	r3, put_sprite_16_aligned.loop
  743=>x"C005",	-- 1100000000000101  li	r5, 0
  744=>x"E383",	-- 1110001110000011  ba	-, r6
  745=>x"C07D",	-- 1100000001111101  li	r5, 15
  746=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  747=>x"6600",	-- 0110011000000000  shr	r0, r0, 3
  748=>x"BBE8",	-- 1011101111101000  brieq	r5, put_sprite_16_aligned
  749=>x"062D",	-- 0000011000101101  dec	r5, r5
  750=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  751=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  752=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  753=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  754=>x"063F",	-- 0000011000111111  dec	r7, r7
  755=>x"D23B",	-- 1101001000111011  sw	r3, r7
  756=>x"0412",	-- 0000010000010010  inc	r2, r2
  757=>x"D011",	-- 1101000000010001  lw	r1, r2
  758=>x"CFF8",	-- 1100111111111000  li	r0, -1
  759=>x"3D40",	-- 0011110101000000  rsr	r0, r0, r5
  760=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  761=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  762=>x"D023",	-- 1101000000100011  lw	r3, r4
  763=>x"2600",	-- 0010011000000000  not	r0, r0
  764=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  765=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  766=>x"E421",	-- 1110010000100001  exw	r1, r4
  767=>x"0424",	-- 0000010000100100  inc	r4, r4
  768=>x"D011",	-- 1101000000010001  lw	r1, r2
  769=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  770=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  771=>x"D023",	-- 1101000000100011  lw	r3, r4
  772=>x"2600",	-- 0010011000000000  not	r0, r0
  773=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  774=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  775=>x"E421",	-- 1110010000100001  exw	r1, r4
  776=>x"0412",	-- 0000010000010010  inc	r2, r2
  777=>x"C098",	-- 1100000010011000  li	r0, 19
  778=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  779=>x"D03B",	-- 1101000000111011  lw	r3, r7
  780=>x"043F",	-- 0000010000111111  inc	r7, r7
  781=>x"061B",	-- 0000011000011011  dec	r3, r3
  782=>x"B91C",	-- 1011100100011100  brine	r3, put_sprite_16.loop
  783=>x"C005",	-- 1100000000000101  li	r5, 0
  784=>x"E383",	-- 1110001110000011  ba	-, r6
  785=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  786=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  787=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  788=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  789=>x"C005",	-- 1100000000000101  li	r5, 0
  790=>x"D020",	-- 1101000000100000  lw	r0, r4
  791=>x"D011",	-- 1101000000010001  lw	r1, r2
  792=>x"0412",	-- 0000010000010010  inc	r2, r2
  793=>x"2040",	-- 0010000001000000  and	r0, r0, r1
  794=>x"D011",	-- 1101000000010001  lw	r1, r2
  795=>x"2240",	-- 0010001001000000  or	r0, r0, r1
  796=>x"E420",	-- 1110010000100000  exw	r0, r4
  797=>x"0612",	-- 0000011000010010  dec	r2, r2
  798=>x"D011",	-- 1101000000010001  lw	r1, r2
  799=>x"2609",	-- 0010011000001001  not	r1, r1
  800=>x"0412",	-- 0000010000010010  inc	r2, r2
  801=>x"2040",	-- 0010000001000000  and	r0, r0, r1
  802=>x"222D",	-- 0010001000101101  or	r5, r5, r0
  803=>x"0412",	-- 0000010000010010  inc	r2, r2
  804=>x"C0A0",	-- 1100000010100000  li	r0, 20
  805=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  806=>x"061B",	-- 0000011000011011  dec	r3, r3
  807=>x"AE5C",	-- 1010111001011100  brine	r3, put_sprite_16_aligned.loop
  808=>x"E383",	-- 1110001110000011  ba	-, r6
  809=>x"C07D",	-- 1100000001111101  li	r5, 15
  810=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  811=>x"6600",	-- 0110011000000000  shr	r0, r0, 3
  812=>x"B968",	-- 1011100101101000  brieq	r5, put_sprite_16_masked_aligned
  813=>x"062D",	-- 0000011000101101  dec	r5, r5
  814=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  815=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  816=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  817=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  818=>x"063F",	-- 0000011000111111  dec	r7, r7
  819=>x"D23E",	-- 1101001000111110  sw	r6, r7
  820=>x"102E",	-- 0001000000101110  mova	r6, r5
  821=>x"C005",	-- 1100000000000101  li	r5, 0
  822=>x"063F",	-- 0000011000111111  dec	r7, r7
  823=>x"D23B",	-- 1101001000111011  sw	r3, r7
  824=>x"063F",	-- 0000011000111111  dec	r7, r7
  825=>x"D23D",	-- 1101001000111101  sw	r5, r7
  826=>x"D010",	-- 1101000000010000  lw	r0, r2
  827=>x"3980",	-- 0011100110000000  rrr	r0, r0, r6
  828=>x"0412",	-- 0000010000010010  inc	r2, r2
  829=>x"D011",	-- 1101000000010001  lw	r1, r2
  830=>x"3989",	-- 0011100110001001  rrr	r1, r1, r6
  831=>x"CFFD",	-- 1100111111111101  li	r5, -1
  832=>x"3DAD",	-- 0011110110101101  rsr	r5, r5, r6
  833=>x"2149",	-- 0010000101001001  and	r1, r1, r5
  834=>x"D023",	-- 1101000000100011  lw	r3, r4
  835=>x"262D",	-- 0010011000101101  not	r5, r5
  836=>x"222D",	-- 0010001000101101  or	r5, r5, r0
  837=>x"215B",	-- 0010000101011011  and	r3, r3, r5
  838=>x"225B",	-- 0010001001011011  or	r3, r3, r1
  839=>x"E423",	-- 1110010000100011  exw	r3, r4
  840=>x"262D",	-- 0010011000101101  not	r5, r5
  841=>x"215B",	-- 0010000101011011  and	r3, r3, r5
  842=>x"D03D",	-- 1101000000111101  lw	r5, r7
  843=>x"043F",	-- 0000010000111111  inc	r7, r7
  844=>x"22ED",	-- 0010001011101101  or	r5, r5, r3
  845=>x"0424",	-- 0000010000100100  inc	r4, r4
  846=>x"063F",	-- 0000011000111111  dec	r7, r7
  847=>x"D23D",	-- 1101001000111101  sw	r5, r7
  848=>x"D011",	-- 1101000000010001  lw	r1, r2
  849=>x"3989",	-- 0011100110001001  rrr	r1, r1, r6
  850=>x"CFFD",	-- 1100111111111101  li	r5, -1
  851=>x"3DAD",	-- 0011110110101101  rsr	r5, r5, r6
  852=>x"262D",	-- 0010011000101101  not	r5, r5
  853=>x"2149",	-- 0010000101001001  and	r1, r1, r5
  854=>x"D023",	-- 1101000000100011  lw	r3, r4
  855=>x"262D",	-- 0010011000101101  not	r5, r5
  856=>x"222D",	-- 0010001000101101  or	r5, r5, r0
  857=>x"215B",	-- 0010000101011011  and	r3, r3, r5
  858=>x"225B",	-- 0010001001011011  or	r3, r3, r1
  859=>x"E423",	-- 1110010000100011  exw	r3, r4
  860=>x"262D",	-- 0010011000101101  not	r5, r5
  861=>x"215B",	-- 0010000101011011  and	r3, r3, r5
  862=>x"D03D",	-- 1101000000111101  lw	r5, r7
  863=>x"043F",	-- 0000010000111111  inc	r7, r7
  864=>x"22ED",	-- 0010001011101101  or	r5, r5, r3
  865=>x"0412",	-- 0000010000010010  inc	r2, r2
  866=>x"C098",	-- 1100000010011000  li	r0, 19
  867=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  868=>x"D03B",	-- 1101000000111011  lw	r3, r7
  869=>x"043F",	-- 0000010000111111  inc	r7, r7
  870=>x"061B",	-- 0000011000011011  dec	r3, r3
  871=>x"B3DC",	-- 1011001111011100  brine	r3, put_sprite_16_masked.loop
  872=>x"D03E",	-- 1101000000111110  lw	r6, r7
  873=>x"043F",	-- 0000010000111111  inc	r7, r7
  874=>x"E383",	-- 1110001110000011  ba	-, r6
  875=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  876=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  877=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  878=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  879=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  880=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  881=>x"C0A5",	-- 1100000010100101  li	r5, 20
  882=>x"8404",	-- 1000010000000100  brine	r0, put_sprite_8_aligned.loop1
  883=>x"D010",	-- 1101000000010000  lw	r0, r2
  884=>x"D021",	-- 1101000000100001  lw	r1, r4
  885=>x"1A41",	-- 0001101001000001  mixhl	r1, r0, r1
  886=>x"D221",	-- 1101001000100001  sw	r1, r4
  887=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  888=>x"061B",	-- 0000011000011011  dec	r3, r3
  889=>x"E398",	-- 1110001110011000  baeq	r3, r6
  890=>x"D021",	-- 1101000000100001  lw	r1, r4
  891=>x"1E41",	-- 0001111001000001  mixll	r1, r0, r1
  892=>x"D221",	-- 1101001000100001  sw	r1, r4
  893=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  894=>x"0412",	-- 0000010000010010  inc	r2, r2
  895=>x"061B",	-- 0000011000011011  dec	r3, r3
  896=>x"E398",	-- 1110001110011000  baeq	r3, r6
  897=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop0
  898=>x"D010",	-- 1101000000010000  lw	r0, r2
  899=>x"D021",	-- 1101000000100001  lw	r1, r4
  900=>x"1809",	-- 0001100000001001  mixhh	r1, r1, r0
  901=>x"D221",	-- 1101001000100001  sw	r1, r4
  902=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  903=>x"061B",	-- 0000011000011011  dec	r3, r3
  904=>x"E398",	-- 1110001110011000  baeq	r3, r6
  905=>x"D021",	-- 1101000000100001  lw	r1, r4
  906=>x"1A09",	-- 0001101000001001  mixhl	r1, r1, r0
  907=>x"D221",	-- 1101001000100001  sw	r1, r4
  908=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  909=>x"0412",	-- 0000010000010010  inc	r2, r2
  910=>x"061B",	-- 0000011000011011  dec	r3, r3
  911=>x"E398",	-- 1110001110011000  baeq	r3, r6
  912=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop1
  913=>x"C03D",	-- 1100000000111101  li	r5, 7
  914=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  915=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  916=>x"B5E8",	-- 1011010111101000  brieq	r5, put_sprite_8_aligned
  917=>x"062D",	-- 0000011000101101  dec	r5, r5
  918=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  919=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  920=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  921=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  922=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  923=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  924=>x"8A04",	-- 1000101000000100  brine	r0, put_sprite_8.loop1
  925=>x"D010",	-- 1101000000010000  lw	r0, r2
  926=>x"063F",	-- 0000011000111111  dec	r7, r7
  927=>x"D23A",	-- 1101001000111010  sw	r2, r7
  928=>x"C802",	-- 1100100000000010  li	r2, 0x100
  929=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  930=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  931=>x"D021",	-- 1101000000100001  lw	r1, r4
  932=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  933=>x"2612",	-- 0010011000010010  not	r2, r2
  934=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  935=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  936=>x"D221",	-- 1101001000100001  sw	r1, r4
  937=>x"C0A1",	-- 1100000010100001  li	r1, 20
  938=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  939=>x"D03A",	-- 1101000000111010  lw	r2, r7
  940=>x"043F",	-- 0000010000111111  inc	r7, r7
  941=>x"061B",	-- 0000011000011011  dec	r3, r3
  942=>x"E398",	-- 1110001110011000  baeq	r3, r6
  943=>x"D010",	-- 1101000000010000  lw	r0, r2
  944=>x"063F",	-- 0000011000111111  dec	r7, r7
  945=>x"D23A",	-- 1101001000111010  sw	r2, r7
  946=>x"1E00",	-- 0001111000000000  mixll	r0, r0, r0
  947=>x"C802",	-- 1100100000000010  li	r2, 0x100
  948=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  949=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  950=>x"D021",	-- 1101000000100001  lw	r1, r4
  951=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  952=>x"2612",	-- 0010011000010010  not	r2, r2
  953=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  954=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  955=>x"D221",	-- 1101001000100001  sw	r1, r4
  956=>x"C0A1",	-- 1100000010100001  li	r1, 20
  957=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  958=>x"D03A",	-- 1101000000111010  lw	r2, r7
  959=>x"043F",	-- 0000010000111111  inc	r7, r7
  960=>x"0412",	-- 0000010000010010  inc	r2, r2
  961=>x"061B",	-- 0000011000011011  dec	r3, r3
  962=>x"E398",	-- 1110001110011000  baeq	r3, r6
  963=>x"B683",	-- 1011011010000011  bri	-, put_sprite_8.loop0
  964=>x"D010",	-- 1101000000010000  lw	r0, r2
  965=>x"063F",	-- 0000011000111111  dec	r7, r7
  966=>x"D23A",	-- 1101001000111010  sw	r2, r7
  967=>x"063F",	-- 0000011000111111  dec	r7, r7
  968=>x"D23B",	-- 1101001000111011  sw	r3, r7
  969=>x"C802",	-- 1100100000000010  li	r2, 0x100
  970=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  971=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  972=>x"2080",	-- 0010000010000000  and	r0, r0, r2
  973=>x"D021",	-- 1101000000100001  lw	r1, r4
  974=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
  975=>x"261B",	-- 0010011000011011  not	r3, r3
  976=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  977=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
  978=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  979=>x"D221",	-- 1101001000100001  sw	r1, r4
  980=>x"0424",	-- 0000010000100100  inc	r4, r4
  981=>x"D021",	-- 1101000000100001  lw	r1, r4
  982=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  983=>x"261B",	-- 0010011000011011  not	r3, r3
  984=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  985=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
  986=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  987=>x"D221",	-- 1101001000100001  sw	r1, r4
  988=>x"C099",	-- 1100000010011001  li	r1, 19
  989=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  990=>x"D03B",	-- 1101000000111011  lw	r3, r7
  991=>x"043F",	-- 0000010000111111  inc	r7, r7
  992=>x"D03A",	-- 1101000000111010  lw	r2, r7
  993=>x"043F",	-- 0000010000111111  inc	r7, r7
  994=>x"061B",	-- 0000011000011011  dec	r3, r3
  995=>x"E398",	-- 1110001110011000  baeq	r3, r6
  996=>x"D010",	-- 1101000000010000  lw	r0, r2
  997=>x"4E00",	-- 0100111000000000  shl	r0, r0, 7
  998=>x"063F",	-- 0000011000111111  dec	r7, r7
  999=>x"D23A",	-- 1101001000111010  sw	r2, r7
 1000=>x"063F",	-- 0000011000111111  dec	r7, r7
 1001=>x"D23B",	-- 1101001000111011  sw	r3, r7
 1002=>x"C802",	-- 1100100000000010  li	r2, 0x100
 1003=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
 1004=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
 1005=>x"2080",	-- 0010000010000000  and	r0, r0, r2
 1006=>x"D021",	-- 1101000000100001  lw	r1, r4
 1007=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
 1008=>x"261B",	-- 0010011000011011  not	r3, r3
 1009=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
 1010=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
 1011=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
 1012=>x"D221",	-- 1101001000100001  sw	r1, r4
 1013=>x"0424",	-- 0000010000100100  inc	r4, r4
 1014=>x"D021",	-- 1101000000100001  lw	r1, r4
 1015=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
 1016=>x"261B",	-- 0010011000011011  not	r3, r3
 1017=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
 1018=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
 1019=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
 1020=>x"D221",	-- 1101001000100001  sw	r1, r4
 1021=>x"C099",	-- 1100000010011001  li	r1, 19
 1022=>x"0864",	-- 0000100001100100  add	r4, r4, r1
 1023=>x"D03B",	-- 1101000000111011  lw	r3, r7
 1024=>x"043F",	-- 0000010000111111  inc	r7, r7
 1025=>x"D03A",	-- 1101000000111010  lw	r2, r7
 1026=>x"043F",	-- 0000010000111111  inc	r7, r7
 1027=>x"0412",	-- 0000010000010010  inc	r2, r2
 1028=>x"061B",	-- 0000011000011011  dec	r3, r3
 1029=>x"E398",	-- 1110001110011000  baeq	r3, r6
 1030=>x"AF83",	-- 1010111110000011  bri	-, put_sprite_8.loop1
    others => x"0000"
    );
begin
  process(CLK)
  begin
    if (CLK'event AND CLK='1') then
      D <= m(to_integer(unsigned(AD)));
    end if;
  end process;
end Behavioral;
