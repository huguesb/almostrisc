----------------------------------------------------------------------------------
--
-- File retrieved, on 07/02/2010, from :
-- http://sebastien-viardot.imag.fr/Enseignements/Archi1A2s/sources/ROMPROG.vhd
--
-- Slightly altered to get rid of vendor-specific packages and adjust formatting
-- Now auto-filled by asrom script
--
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROMPROG is
  Port ( AD : in  STD_LOGIC_VECTOR (12 downto 0);
         D : out  STD_LOGIC_VECTOR (15 downto 0);
         CLK : in STD_LOGIC);
end ROMPROG;

architecture Behavioral of ROMPROG is
  constant low_address: natural := 0;
  constant high_address: natural := 8192;
  subtype octet is std_logic_vector( 15 downto 0 );
  type zone_memoire is
    array (natural range low_address to high_address-1) of octet;
  constant m: zone_memoire:= (
    0=>x"FFF7",	-- 1111111111110111  liw	r7, IRQ_mask
    1=>x"2000",	-- 0010000000000000  
    2=>x"F8C0",	-- 1111100011000000  bai	-, os_init
    3=>x"0100",	-- 0000000100000000  
   16=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_ack
   17=>x"2002",	-- 0010000000000010  
   18=>x"D001",	-- 1101000000000001  lw	r1, r0
   19=>x"F54A",	-- 1111010101001010  bspl	r2, r1, 5
   20=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_error
   21=>x"0050",	-- 0000000001010000  
   22=>x"F4CA",	-- 1111010011001010  bspl	r2, r1, 3
   23=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_kbd
   24=>x"0060",	-- 0000000001100000  
   25=>x"F40A",	-- 1111010000001010  bspl	r2, r1, 0
   26=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_tmr
   27=>x"0040",	-- 0000000001000000  
   28=>x"D201",	-- 1101001000000001  sw	r1, r0
   29=>x"FFFE",	-- 1111111111111110  reti
   64=>x"263F",	-- 0010011000111111  not r7, r7
   65=>x"D7C0",	-- 1101011111000000  out	r7
   66=>x"E383",	-- 1110001110000011  ba	-, r6
   80=>x"25FF",	-- 0010010111111111  xor	r7, r7, r7
   81=>x"D7C0",	-- 1101011111000000  out	r7
   82=>x"E383",	-- 1110001110000011  ba	-, r6
   96=>x"FFF2",	-- 1111111111110010  liw	r2, PS2_rx
   97=>x"2004",	-- 0010000000000100  
   98=>x"D012",	-- 1101000000010010  lw	r2, r2
   99=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map + 8
  100=>x"1808",	-- 0001100000001000  
  101=>x"D01B",	-- 1101000000011011  lw	r3, r3
  102=>x"1EBF",	-- 0001111010111111  mixll	r7, r7, r2
  103=>x"C784",	-- 1100011110000100  li	r4, 0xF0
  104=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  105=>x"8B20",	-- 1000101100100000  brieq	r4, int_kbd.release
  106=>x"C704",	-- 1100011100000100  li	r4, 0xE0
  107=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  108=>x"88E0",	-- 1000100011100000  brieq	r4, int_kbd.extended
  109=>x"FFF5",	-- 1111111111110101  liw	r5, paper_keys - 1
  110=>x"16BF",	-- 0001011010111111  
  111=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  112=>x"80E0",	-- 1000000011100000  brieq	r4, $+3
  113=>x"FFF5",	-- 1111111111110101  liw	r5, paper_keys + 10 - 1
  114=>x"16C9",	-- 0001011011001001  
  115=>x"042D",	-- 0000010000101101  inc	r5, r5
  116=>x"D02C",	-- 1101000000101100  lw	r4, r5
  117=>x"8560",	-- 1000010101100000  brieq	r4, scan_code_mismatch
  118=>x"6E24",	-- 0110111000100100  shr	r4, r4, 7
  119=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  120=>x"BEE4",	-- 1011111011100100  brine	r4, scan_code_loop
  121=>x"D02A",	-- 1101000000101010  lw	r2, r5
  122=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  123=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  124=>x"741B",	-- 0111010000011011  shr	r3, r3, 10
  125=>x"C00D",	-- 1100000000001101  li	r5, 1
  126=>x"0612",	-- 0000011000010010  dec	r2, r2
  127=>x"3AAA",	-- 0011101010101010  rrl	r2, r5, r2
  128=>x"FFF5",	-- 1111111111110101  liw	r5, key_press_map
  129=>x"1800",	-- 0001100000000000  
  130=>x"08ED",	-- 0000100011101101  add	r5, r5, r3
  131=>x"D02B",	-- 1101000000101011  lw	r3, r5
  132=>x"80E4",	-- 1000000011100100  brine	r4, scan_code_release
  133=>x"229B",	-- 0010001010011011  or	r3, r3, r2
  134=>x"80C3",	-- 1000000011000011  bri	-, scan_code_notify
  135=>x"2612",	-- 0010011000010010  not	r2, r2
  136=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  137=>x"D22B",	-- 1101001000101011  sw	r3, r5
  138=>x"C003",	-- 1100000000000011  li	r3, 0
  139=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  140=>x"1808",	-- 0001100000001000  
  141=>x"D223",	-- 1101001000100011  sw	r3, r4
  142=>x"E383",	-- 1110001110000011  ba	-, r6
  143=>x"C014",	-- 1100000000010100  li	r4, 2
  144=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  145=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  146=>x"1808",	-- 0001100000001000  
  147=>x"D223",	-- 1101001000100011  sw	r3, r4
  148=>x"E383",	-- 1110001110000011  ba	-, r6
  149=>x"C00C",	-- 1100000000001100  li	r4, 1
  150=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  151=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  152=>x"1808",	-- 0001100000001000  
  153=>x"D223",	-- 1101001000100011  sw	r3, r4
  154=>x"E383",	-- 1110001110000011  ba	-, r6
  256=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_mask
  257=>x"2000",	-- 0010000000000000  
  258=>x"C0C9",	-- 1100000011001001  li	r1, 0x19
  259=>x"D201",	-- 1101001000000001  sw	r1, r0
  260=>x"0400",	-- 0000010000000000  inc	r0, r0
  261=>x"CFF9",	-- 1100111111111001  li	r1, -1
  262=>x"D201",	-- 1101001000000001  sw	r1, r0
  263=>x"C03A",	-- 1100000000111010  li	r2, 7
  264=>x"0880",	-- 0000100010000000  add	r0, r0, r2
  265=>x"C0EA",	-- 1100000011101010  li	r2, 0x1D
  266=>x"D202",	-- 1101001000000010  sw	r2, r0
  267=>x"0400",	-- 0000010000000000  inc	r0, r0
  268=>x"C07A",	-- 1100000001111010  li	r2, 15
  269=>x"D202",	-- 1101001000000010  sw	r2, r0
  270=>x"FFF0",	-- 1111111111110000  liw	r0, key_press_map
  271=>x"1800",	-- 0001100000000000  
  272=>x"C001",	-- 1100000000000001  li	r1, 0
  273=>x"C042",	-- 1100000001000010  li	r2, 8
  274=>x"D201",	-- 1101001000000001  sw	r1, r0
  275=>x"0400",	-- 0000010000000000  inc	r0, r0
  276=>x"0612",	-- 0000011000010010  dec	r2, r2
  277=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  278=>x"C0F3",	-- 1100000011110011  li	r3, 30
  279=>x"CFFA",	-- 1100111111111010  li	r2, -1
  280=>x"D21A",	-- 1101001000011010  sw	r2, r3
  281=>x"8083",	-- 1000000010000011  bri	-, PaperGameStart
  282=>x"8003",	-- 1000000000000011  bri	-, PaperMenuLoop
  283=>x"FFF0",	-- 1111111111110000  liw	r0, paper_dir
  284=>x"1730",	-- 0001011100110000  
  285=>x"C001",	-- 1100000000000001  li	r1, 0
  286=>x"D201",	-- 1101001000000001  sw	r1, r0
  287=>x"0400",	-- 0000010000000000  inc	r0, r0
  288=>x"C4C1",	-- 1100010011000001  li	r1, 152
  289=>x"D201",	-- 1101001000000001  sw	r1, r0
  290=>x"0400",	-- 0000010000000000  inc	r0, r0
  291=>x"C001",	-- 1100000000000001  li	r1, 0
  292=>x"D201",	-- 1101001000000001  sw	r1, r0
  293=>x"0400",	-- 0000010000000000  inc	r0, r0
  294=>x"C401",	-- 1100010000000001  li	r1, 128
  295=>x"D201",	-- 1101001000000001  sw	r1, r0
  296=>x"0400",	-- 0000010000000000  inc	r0, r0
  297=>x"C001",	-- 1100000000000001  li	r1, 0
  298=>x"D201",	-- 1101001000000001  sw	r1, r0
  299=>x"0400",	-- 0000010000000000  inc	r0, r0
  300=>x"C0A1",	-- 1100000010100001  li	r1, 20
  301=>x"D201",	-- 1101001000000001  sw	r1, r0
  302=>x"0400",	-- 0000010000000000  inc	r0, r0
  303=>x"C029",	-- 1100000000101001  li	r1, 5
  304=>x"D201",	-- 1101001000000001  sw	r1, r0
  305=>x"0400",	-- 0000010000000000  inc	r0, r0
  306=>x"C000",	-- 1100000000000000  li	r0, 0
  307=>x"CFF9",	-- 1100111111111001  li	r1, -1
  308=>x"C0A2",	-- 1100000010100010  li	r2, 20
  309=>x"D201",	-- 1101001000000001  sw	r1, r0
  310=>x"0400",	-- 0000010000000000  inc	r0, r0
  311=>x"0612",	-- 0000011000010010  dec	r2, r2
  312=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  313=>x"C001",	-- 1100000000000001  li	r1, 0
  314=>x"FFF2",	-- 1111111111110010  liw	r2, 18*20
  315=>x"0168",	-- 0000000101101000  
  316=>x"D201",	-- 1101001000000001  sw	r1, r0
  317=>x"0400",	-- 0000010000000000  inc	r0, r0
  318=>x"0612",	-- 0000011000010010  dec	r2, r2
  319=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  320=>x"CFF9",	-- 1100111111111001  li	r1, -1
  321=>x"C0A2",	-- 1100000010100010  li	r2, 20
  322=>x"D201",	-- 1101001000000001  sw	r1, r0
  323=>x"0400",	-- 0000010000000000  inc	r0, r0
  324=>x"0612",	-- 0000011000010010  dec	r2, r2
  325=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  326=>x"C020",	-- 1100000000100000  li	r0, 4
  327=>x"C029",	-- 1100000000101001  li	r1, 5
  328=>x"FFF2",	-- 1111111111110010  liw	r2, paper_title
  329=>x"1738",	-- 0001011100111000  
  330=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  331=>x"01CB",	-- 0000000111001011  
  332=>x"C790",	-- 1100011110010000  li	r0, 242
  333=>x"C009",	-- 1100000000001001  li	r1, 1
  334=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud
  335=>x"1720",	-- 0001011100100000  
  336=>x"C043",	-- 1100000001000011  li	r3, 8
  337=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  338=>x"0256",	-- 0000001001010110  
  339=>x"C118",	-- 1100000100011000  li	r0, 35
  340=>x"C009",	-- 1100000000001001  li	r1, 1
  341=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  342=>x"173E",	-- 0001011100111110  
  343=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  344=>x"01CB",	-- 0000000111001011  
  345=>x"C790",	-- 1100011110010000  li	r0, 242
  346=>x"C051",	-- 1100000001010001  li	r1, 10
  347=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud + 4
  348=>x"1724",	-- 0001011100100100  
  349=>x"C043",	-- 1100000001000011  li	r3, 8
  350=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  351=>x"0256",	-- 0000001001010110  
  352=>x"C118",	-- 1100000100011000  li	r0, 35
  353=>x"C051",	-- 1100000001010001  li	r1, 10
  354=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  355=>x"173E",	-- 0001011100111110  
  356=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  357=>x"01CB",	-- 0000000111001011  
  358=>x"FFF0",	-- 1111111111110000  liw	r0, 20*20
  359=>x"0190",	-- 0000000110010000  
  360=>x"C001",	-- 1100000000000001  li	r1, 0
  361=>x"FFF2",	-- 1111111111110010  liw	r2, 220*20
  362=>x"1130",	-- 0001000100110000  
  363=>x"D201",	-- 1101001000000001  sw	r1, r0
  364=>x"0400",	-- 0000010000000000  inc	r0, r0
  365=>x"0612",	-- 0000011000010010  dec	r2, r2
  366=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  367=>x"FFF3",	-- 1111111111110011  liw	r3, paper_dir
  368=>x"1730",	-- 0001011100110000  
  369=>x"D01C",	-- 1101000000011100  lw	r4, r3
  370=>x"041B",	-- 0000010000011011  inc	r3, r3
  371=>x"D018",	-- 1101000000011000  lw	r0, r3
  372=>x"FFF2",	-- 1111111111110010  liw	r2, paper_sprites
  373=>x"16D0",	-- 0001011011010000  
  374=>x"4624",	-- 0100011000100100  shl	r4, r4, 3
  375=>x"0912",	-- 0000100100010010  add	r2, r2, r4
  376=>x"C161",	-- 1100000101100001  li	r1, 44
  377=>x"C083",	-- 1100000010000011  li	r3, 16
  378=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_16
  379=>x"0206",	-- 0000001000000110  
  380=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  381=>x"1800",	-- 0001100000000000  
  382=>x"D01B",	-- 1101000000011011  lw	r3, r3
  383=>x"BF58",	-- 1011111101011000  brieq	r3, PaperGameLoop
  384=>x"F7DC",	-- 1111011111011100  bspl	r4, r3, 15
  385=>x"86A4",	-- 1000011010100100  brine	r4, PaperGameQuit
  386=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  387=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveUp
  388=>x"F49C",	-- 1111010010011100  bspl	r4, r3, 2
  389=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveDOWN
  390=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  391=>x"8260",	-- 1000001001100000  brieq	r4, PaperNoMoveLEFT
  392=>x"FFF2",	-- 1111111111110010  liw	r2, paper_dir
  393=>x"1730",	-- 0001011100110000  
  394=>x"C010",	-- 1100000000010000  li	r0, 2
  395=>x"D210",	-- 1101001000010000  sw	r0, r2
  396=>x"0412",	-- 0000010000010010  inc	r2, r2
  397=>x"D010",	-- 1101000000010000  lw	r0, r2
  398=>x"0600",	-- 0000011000000000  dec	r0, r0
  399=>x"D210",	-- 1101001000010000  sw	r0, r2
  400=>x"F4DC",	-- 1111010011011100  bspl	r4, r3, 3
  401=>x"8260",	-- 1000001001100000  brieq	r4, PaperNoMoveRIGHT
  402=>x"FFF2",	-- 1111111111110010  liw	r2, paper_dir
  403=>x"1730",	-- 0001011100110000  
  404=>x"C008",	-- 1100000000001000  li	r0, 1
  405=>x"D210",	-- 1101001000010000  sw	r0, r2
  406=>x"0412",	-- 0000010000010010  inc	r2, r2
  407=>x"D010",	-- 1101000000010000  lw	r0, r2
  408=>x"0400",	-- 0000010000000000  inc	r0, r0
  409=>x"D210",	-- 1101001000010000  sw	r0, r2
  410=>x"B303",	-- 1011001100000011  bri	-, PaperGameRedrawContent
  411=>x"FFFF",	-- 1111111111111111  reset
  412=>x"C750",	-- 1100011101010000  li	r0, 234
  413=>x"C1C2",	-- 1100000111000010  li	r2, 56
  414=>x"FAC6",	-- 1111101011000110  bail	-, r6, div_16_16
  415=>x"01B4",	-- 0000000110110100  
  416=>x"C448",	-- 1100010001001000  li	r0, 137
  417=>x"C472",	-- 1100010001110010  li	r2, 142
  418=>x"FAC6",	-- 1111101011000110  bail	-, r6, mult_16_16
  419=>x"01A8",	-- 0000000110101000  
  420=>x"C03A",	-- 1100000000111010  li r2, 7
  421=>x"FAC6",	-- 1111101011000110  bail	-, r6, fact_16
  422=>x"01BF",	-- 0000000110111111  
  423=>x"FFFF",	-- 1111111111111111  reset
  424=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  425=>x"2524",	-- 0010010100100100  xor	r4, r4, r4
  426=>x"C085",	-- 1100000010000101  li	r5, 16
  427=>x"0849",	-- 0000100001001001  add	r1, r1, r1
  428=>x"0C00",	-- 0000110000000000  adc	r0, r0, r0
  429=>x"0EDB",	-- 0000111011011011  sbc	r3, r3, r3
  430=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  431=>x"08C9",	-- 0000100011001001  add	r1, r1, r3
  432=>x"0D00",	-- 0000110100000000  adc	r0, r0, r4
  433=>x"062D",	-- 0000011000101101  dec	r5, r5
  434=>x"BE6C",	-- 1011111001101100  brine	r5, mult_16_16.loop
  435=>x"E383",	-- 1110001110000011  ba	-, r6
  436=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  437=>x"C084",	-- 1100000010000100  li	r4, 16
  438=>x"0800",	-- 0000100000000000  add	r0, r0, r0
  439=>x"0C49",	-- 0000110001001001  adc	r1, r1, r1
  440=>x"0A8B",	-- 0000101010001011  sub	r3, r1, r2
  441=>x"80DD",	-- 1000000011011101  brilt	r3, div_16_16.skip
  442=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  443=>x"0400",	-- 0000010000000000  inc	r0, r0
  444=>x"0624",	-- 0000011000100100  dec	r4, r4
  445=>x"BE64",	-- 1011111001100100  brine	r4, div_16_16.loop
  446=>x"E383",	-- 1110001110000011  ba	-, r6
  447=>x"2400",	-- 0010010000000000  xor	r0, r0, r0
  448=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  449=>x"8250",	-- 1000001001010000  brieq	r2, fact_16.end
  450=>x"0409",	-- 0000010000001001  inc	r1, r1
  451=>x"1008",	-- 0001000000001000  mova	r0, r1
  452=>x"FAC6",	-- 1111101011000110  bail	-, r6, mult_16_16
  453=>x"01A8",	-- 0000000110101000  
  454=>x"8104",	-- 1000000100000100  brine	r0, fact_16.overflow
  455=>x"01A8",	-- 0000000110101000  
  456=>x"0612",	-- 0000011000010010  dec	r2, r2
  457=>x"BE94",	-- 1011111010010100  brine	r2, fact_16.loop
  458=>x"E383",	-- 1110001110000011  ba	-, r6
  459=>x"063F",	-- 0000011000111111  dec	r7, r7
  460=>x"D23E",	-- 1101001000111110  sw	r6, r7
  461=>x"D013",	-- 1101000000010011  lw	r3, r2
  462=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  463=>x"84D8",	-- 1000010011011000  brieq	r3, puts.end
  464=>x"063F",	-- 0000011000111111  dec	r7, r7
  465=>x"D23A",	-- 1101001000111010  sw	r2, r7
  466=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  467=>x"01E5",	-- 0000000111100101  
  468=>x"D03A",	-- 1101000000111010  lw	r2, r7
  469=>x"043F",	-- 0000010000111111  inc	r7, r7
  470=>x"D013",	-- 1101000000010011  lw	r3, r2
  471=>x"4E1B",	-- 0100111000011011  shl	r3, r3, 7
  472=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  473=>x"8258",	-- 1000001001011000  brieq	r3, puts.end
  474=>x"063F",	-- 0000011000111111  dec	r7, r7
  475=>x"D23A",	-- 1101001000111010  sw	r2, r7
  476=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  477=>x"01E5",	-- 0000000111100101  
  478=>x"D03A",	-- 1101000000111010  lw	r2, r7
  479=>x"043F",	-- 0000010000111111  inc	r7, r7
  480=>x"0412",	-- 0000010000010010  inc	r2, r2
  481=>x"BB03",	-- 1011101100000011  bri	-, puts.loop
  482=>x"D03E",	-- 1101000000111110  lw	r6, r7
  483=>x"043F",	-- 0000010000111111  inc	r7, r7
  484=>x"E383",	-- 1110001110000011  ba	-, r6
  485=>x"063F",	-- 0000011000111111  dec	r7, r7
  486=>x"D23E",	-- 1101001000111110  sw	r6, r7
  487=>x"063F",	-- 0000011000111111  dec	r7, r7
  488=>x"D238",	-- 1101001000111000  sw	r0, r7
  489=>x"063F",	-- 0000011000111111  dec	r7, r7
  490=>x"D239",	-- 1101001000111001  sw	r1, r7
  491=>x"FFF2",	-- 1111111111110010  liw	r2, font_map
  492=>x"12C0",	-- 0001001011000000  
  493=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  494=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  495=>x"C043",	-- 1100000001000011  li	r3, 8
  496=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  497=>x"0230",	-- 0000001000110000  
  498=>x"D039",	-- 1101000000111001  lw	r1, r7
  499=>x"043F",	-- 0000010000111111  inc	r7, r7
  500=>x"D038",	-- 1101000000111000  lw	r0, r7
  501=>x"043F",	-- 0000010000111111  inc	r7, r7
  502=>x"0400",	-- 0000010000000000  inc	r0, r0
  503=>x"D03E",	-- 1101000000111110  lw	r6, r7
  504=>x"043F",	-- 0000010000111111  inc	r7, r7
  505=>x"E383",	-- 1110001110000011  ba	-, r6
  506=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  507=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  508=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  509=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  510=>x"C0A0",	-- 1100000010100000  li	r0, 20
  511=>x"D011",	-- 1101000000010001  lw	r1, r2
  512=>x"D221",	-- 1101001000100001  sw	r1, r4
  513=>x"0412",	-- 0000010000010010  inc	r2, r2
  514=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  515=>x"061B",	-- 0000011000011011  dec	r3, r3
  516=>x"BEDC",	-- 1011111011011100  brine	r3, put_sprite_16_aligned.loop
  517=>x"E383",	-- 1110001110000011  ba	-, r6
  518=>x"C07D",	-- 1100000001111101  li	r5, 15
  519=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  520=>x"6600",	-- 0110011000000000  shr	r0, r0, 3
  521=>x"BC68",	-- 1011110001101000  brieq	r5, put_sprite_16_aligned
  522=>x"062D",	-- 0000011000101101  dec	r5, r5
  523=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  524=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  525=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  526=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  527=>x"063F",	-- 0000011000111111  dec	r7, r7
  528=>x"D23B",	-- 1101001000111011  sw	r3, r7
  529=>x"D011",	-- 1101000000010001  lw	r1, r2
  530=>x"CFF8",	-- 1100111111111000  li	r0, -1
  531=>x"3D40",	-- 0011110101000000  rsr	r0, r0, r5
  532=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  533=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  534=>x"D023",	-- 1101000000100011  lw	r3, r4
  535=>x"2600",	-- 0010011000000000  not	r0, r0
  536=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  537=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  538=>x"D221",	-- 1101001000100001  sw	r1, r4
  539=>x"0424",	-- 0000010000100100  inc	r4, r4
  540=>x"D011",	-- 1101000000010001  lw	r1, r2
  541=>x"262D",	-- 0010011000101101  not	r5, r5
  542=>x"CFF8",	-- 1100111111111000  li	r0, -1
  543=>x"3F40",	-- 0011111101000000  rsl	r0, r0, r5
  544=>x"3B49",	-- 0011101101001001  rrl	r1, r1, r5
  545=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  546=>x"262D",	-- 0010011000101101  not	r5, r5
  547=>x"D023",	-- 1101000000100011  lw	r3, r4
  548=>x"2600",	-- 0010011000000000  not	r0, r0
  549=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  550=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  551=>x"D221",	-- 1101001000100001  sw	r1, r4
  552=>x"0412",	-- 0000010000010010  inc	r2, r2
  553=>x"C098",	-- 1100000010011000  li	r0, 19
  554=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  555=>x"D03B",	-- 1101000000111011  lw	r3, r7
  556=>x"043F",	-- 0000010000111111  inc	r7, r7
  557=>x"061B",	-- 0000011000011011  dec	r3, r3
  558=>x"B85C",	-- 1011100001011100  brine	r3, put_sprite_16.loop
  559=>x"E383",	-- 1110001110000011  ba	-, r6
  560=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  561=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  562=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  563=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  564=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  565=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  566=>x"C0A5",	-- 1100000010100101  li	r5, 20
  567=>x"8404",	-- 1000010000000100  brine	r0, put_sprite_8_aligned.loop1
  568=>x"D010",	-- 1101000000010000  lw	r0, r2
  569=>x"D021",	-- 1101000000100001  lw	r1, r4
  570=>x"1A41",	-- 0001101001000001  mixhl	r1, r0, r1
  571=>x"D221",	-- 1101001000100001  sw	r1, r4
  572=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  573=>x"061B",	-- 0000011000011011  dec	r3, r3
  574=>x"E398",	-- 1110001110011000  baeq	r3, r6
  575=>x"D021",	-- 1101000000100001  lw	r1, r4
  576=>x"1E41",	-- 0001111001000001  mixll	r1, r0, r1
  577=>x"D221",	-- 1101001000100001  sw	r1, r4
  578=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  579=>x"0412",	-- 0000010000010010  inc	r2, r2
  580=>x"061B",	-- 0000011000011011  dec	r3, r3
  581=>x"E398",	-- 1110001110011000  baeq	r3, r6
  582=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop0
  583=>x"D010",	-- 1101000000010000  lw	r0, r2
  584=>x"D021",	-- 1101000000100001  lw	r1, r4
  585=>x"1809",	-- 0001100000001001  mixhh	r1, r1, r0
  586=>x"D221",	-- 1101001000100001  sw	r1, r4
  587=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  588=>x"061B",	-- 0000011000011011  dec	r3, r3
  589=>x"E398",	-- 1110001110011000  baeq	r3, r6
  590=>x"D021",	-- 1101000000100001  lw	r1, r4
  591=>x"1A09",	-- 0001101000001001  mixhl	r1, r1, r0
  592=>x"D221",	-- 1101001000100001  sw	r1, r4
  593=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  594=>x"0412",	-- 0000010000010010  inc	r2, r2
  595=>x"061B",	-- 0000011000011011  dec	r3, r3
  596=>x"E398",	-- 1110001110011000  baeq	r3, r6
  597=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop1
  598=>x"C03D",	-- 1100000000111101  li	r5, 7
  599=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  600=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  601=>x"B5E8",	-- 1011010111101000  brieq	r5, put_sprite_8_aligned
  602=>x"062D",	-- 0000011000101101  dec	r5, r5
  603=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  604=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  605=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  606=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  607=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  608=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  609=>x"8A04",	-- 1000101000000100  brine	r0, put_sprite_8.loop1
  610=>x"D010",	-- 1101000000010000  lw	r0, r2
  611=>x"063F",	-- 0000011000111111  dec	r7, r7
  612=>x"D23A",	-- 1101001000111010  sw	r2, r7
  613=>x"C802",	-- 1100100000000010  li	r2, 0x100
  614=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  615=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  616=>x"D021",	-- 1101000000100001  lw	r1, r4
  617=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  618=>x"2612",	-- 0010011000010010  not	r2, r2
  619=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  620=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  621=>x"D221",	-- 1101001000100001  sw	r1, r4
  622=>x"C0A1",	-- 1100000010100001  li	r1, 20
  623=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  624=>x"D03A",	-- 1101000000111010  lw	r2, r7
  625=>x"043F",	-- 0000010000111111  inc	r7, r7
  626=>x"061B",	-- 0000011000011011  dec	r3, r3
  627=>x"E398",	-- 1110001110011000  baeq	r3, r6
  628=>x"D010",	-- 1101000000010000  lw	r0, r2
  629=>x"063F",	-- 0000011000111111  dec	r7, r7
  630=>x"D23A",	-- 1101001000111010  sw	r2, r7
  631=>x"1E00",	-- 0001111000000000  mixll	r0, r0, r0
  632=>x"C802",	-- 1100100000000010  li	r2, 0x100
  633=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  634=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  635=>x"D021",	-- 1101000000100001  lw	r1, r4
  636=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  637=>x"2612",	-- 0010011000010010  not	r2, r2
  638=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  639=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  640=>x"D221",	-- 1101001000100001  sw	r1, r4
  641=>x"C0A1",	-- 1100000010100001  li	r1, 20
  642=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  643=>x"D03A",	-- 1101000000111010  lw	r2, r7
  644=>x"043F",	-- 0000010000111111  inc	r7, r7
  645=>x"0412",	-- 0000010000010010  inc	r2, r2
  646=>x"061B",	-- 0000011000011011  dec	r3, r3
  647=>x"E398",	-- 1110001110011000  baeq	r3, r6
  648=>x"B683",	-- 1011011010000011  bri	-, put_sprite_8.loop0
  649=>x"D010",	-- 1101000000010000  lw	r0, r2
  650=>x"063F",	-- 0000011000111111  dec	r7, r7
  651=>x"D23A",	-- 1101001000111010  sw	r2, r7
  652=>x"063F",	-- 0000011000111111  dec	r7, r7
  653=>x"D23B",	-- 1101001000111011  sw	r3, r7
  654=>x"C802",	-- 1100100000000010  li	r2, 0x100
  655=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  656=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  657=>x"2080",	-- 0010000010000000  and	r0, r0, r2
  658=>x"D021",	-- 1101000000100001  lw	r1, r4
  659=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
  660=>x"261B",	-- 0010011000011011  not	r3, r3
  661=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  662=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
  663=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  664=>x"D221",	-- 1101001000100001  sw	r1, r4
  665=>x"0424",	-- 0000010000100100  inc	r4, r4
  666=>x"D021",	-- 1101000000100001  lw	r1, r4
  667=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  668=>x"261B",	-- 0010011000011011  not	r3, r3
  669=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  670=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
  671=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  672=>x"D221",	-- 1101001000100001  sw	r1, r4
  673=>x"C099",	-- 1100000010011001  li	r1, 19
  674=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  675=>x"D03B",	-- 1101000000111011  lw	r3, r7
  676=>x"043F",	-- 0000010000111111  inc	r7, r7
  677=>x"D03A",	-- 1101000000111010  lw	r2, r7
  678=>x"043F",	-- 0000010000111111  inc	r7, r7
  679=>x"061B",	-- 0000011000011011  dec	r3, r3
  680=>x"E398",	-- 1110001110011000  baeq	r3, r6
  681=>x"D010",	-- 1101000000010000  lw	r0, r2
  682=>x"4E00",	-- 0100111000000000  shl	r0, r0, 7
  683=>x"063F",	-- 0000011000111111  dec	r7, r7
  684=>x"D23A",	-- 1101001000111010  sw	r2, r7
  685=>x"063F",	-- 0000011000111111  dec	r7, r7
  686=>x"D23B",	-- 1101001000111011  sw	r3, r7
  687=>x"C802",	-- 1100100000000010  li	r2, 0x100
  688=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  689=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  690=>x"2080",	-- 0010000010000000  and	r0, r0, r2
  691=>x"D021",	-- 1101000000100001  lw	r1, r4
  692=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
  693=>x"261B",	-- 0010011000011011  not	r3, r3
  694=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  695=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
  696=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  697=>x"D221",	-- 1101001000100001  sw	r1, r4
  698=>x"0424",	-- 0000010000100100  inc	r4, r4
  699=>x"D021",	-- 1101000000100001  lw	r1, r4
  700=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  701=>x"261B",	-- 0010011000011011  not	r3, r3
  702=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  703=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
  704=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  705=>x"D221",	-- 1101001000100001  sw	r1, r4
  706=>x"C099",	-- 1100000010011001  li	r1, 19
  707=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  708=>x"D03B",	-- 1101000000111011  lw	r3, r7
  709=>x"043F",	-- 0000010000111111  inc	r7, r7
  710=>x"D03A",	-- 1101000000111010  lw	r2, r7
  711=>x"043F",	-- 0000010000111111  inc	r7, r7
  712=>x"0412",	-- 0000010000010010  inc	r2, r2
  713=>x"061B",	-- 0000011000011011  dec	r3, r3
  714=>x"E398",	-- 1110001110011000  baeq	r3, r6
  715=>x"AF83",	-- 1010111110000011  bri	-, put_sprite_8.loop1
    others => x"0000"
    );
begin
  process(CLK)
  begin
    if (CLK'event AND CLK='1') then
      D <= m(to_integer(unsigned(AD)));
    end if;
  end process;
end Behavioral;
