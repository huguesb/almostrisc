----------------------------------------------------------------------------------
--
-- File retrieved, on 07/02/2010, from :
-- http://sebastien-viardot.imag.fr/Enseignements/Archi1A2s/sources/ROMPROG.vhd
--
-- Slightly altered to get rid of vendor-specific packages and adjust formatting
--
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROMPROG is
  Port ( AD : in  STD_LOGIC_VECTOR (12 downto 0);
         D : out  STD_LOGIC_VECTOR (15 downto 0);
         CLK : in STD_LOGIC);
end ROMPROG;

architecture Behavioral of ROMPROG is
  constant low_address: natural := 0;
  constant high_address: natural := 8192;
  subtype octet is std_logic_vector( 15 downto 0 );
  type zone_memoire is
    array (natural range low_address to high_address-1) of octet;
  constant m: zone_memoire:= (
0=>x"25FF",     -- 0010010111111111  xor        r7, r7, r7
1=>x"F8C0",     -- 1111100011000000  bai        -, os_init
2=>x"0100",     -- 0000000100000000

16=>x"C100",    -- 1100000100000000  li r0, 0x20
17=>x"4E00",    -- 0100111000000000  shl        r0, r0, 7
18=>x"C012",    -- 1100000000010010  li r2, 2
19=>x"0880",    -- 0000100010000000  add        r0, r0, r2
20=>x"CFF9",    -- 1100111111111001  li r1, -1
21=>x"D201",    -- 1101001000000001  sw r1, r0
22=>x"261B",    -- 0010011000011011  not r3, r3
23=>x"D6C0",    -- 1101011011000000  out        r3
24=>x"FFFE",    -- 1111111111111110  reti

256=>x"FFF0",   -- 1111111111110000  liw        r0, 0x2000
257=>x"2000",   -- 0010000000000000  
258=>x"C009",   -- 1100000000001001  li r1, 1
259=>x"D201",   -- 1101001000000001  sw r1, r0
260=>x"0400",   -- 0000010000000000  inc        r0, r0
261=>x"CFF9",   -- 1100111111111001  li r1, -1
262=>x"D201",   -- 1101001000000001  sw r1, r0
263=>x"C03A",   -- 1100000000111010  li r2, 7
264=>x"0880",   -- 0000100010000000  add        r0, r0, r2
265=>x"C0C2",   -- 1100000011000010  li r2, 0x18
266=>x"D202",   -- 1101001000000010  sw r2, r0
267=>x"0400",   -- 0000010000000000  inc        r0, r0
268=>x"C012",   -- 1100000000010010  li r2, 2
269=>x"D202",   -- 1101001000000010  sw r2, r0

270=>x"FFF0",   -- 1111111111110000  liw        r0, 0x8421
271=>x"8421",   -- 1000010000100001  
272=>x"FFF1",   -- 1111111111110001  liw        r1, 0x1234
273=>x"1234",   -- 0001001000110100  
274=>x"E408",   -- 1110010000001000  exw        r0, r1
275=>x"E408",   -- 1110010000001000  exw        r0, r1
276=>x"1842",   -- 0001100001000010  mixhh      r2, r0, r1
277=>x"1A43",   -- 0001101001000011  mixhl      r3, r0, r1
278=>x"1C44",   -- 0001110001000100  mixlh      r4, r0, r1
279=>x"1E45",   -- 0001111001000101  mixll      r5, r0, r1

280=>x"C750",   -- 1100011101010000  li r0, 234
281=>x"C1C2",   -- 1100000111000010  li r2, 56
282=>x"FAF0",   -- 1111101011110000  bail       -, r6, div_16_16
283=>x"0132",   -- 0000000100110010  
284=>x"FFFF",   -- 1111111111111111  reset

285=>x"C448",   -- 1100010001001000  li r0, 137
286=>x"C472",   -- 1100010001110010  li r2, 142
287=>x"FAF0",   -- 1111101011110000  bail       -, r6, mult_16_16
288=>x"0126",   -- 0000000100100110  
289=>x"FFFF",   -- 1111111111111111  reset

290=>x"C03A",   -- 1100000000111010  li r2, 7
291=>x"FAF0",   -- 1111101011110000  bail       -, r6, fact_16
292=>x"013D",   -- 0000000100111101 
293=>x"FFFF",   -- 1111111111111111  reset

294=>x"2449",   -- 0010010001001001  xor        r1, r1, r1
295=>x"2524",   -- 0010010100100100  xor        r4, r4, r4
296=>x"C085",   -- 1100000010000101  li r5, 16
297=>x"0849",   -- 0000100001001001  add        r1, r1, r1
298=>x"0C00",   -- 0000110000000000  adc        r0, r0, r0
299=>x"0EDB",   -- 0000111011011011  sbc        r3, r3, r3
300=>x"209B",   -- 0010000010011011  and        r3, r3, r2
301=>x"08C9",   -- 0000100011001001  add        r1, r1, r3
302=>x"0D00",   -- 0000110100000000  adc        r0, r0, r4
303=>x"062D",   -- 0000011000101101  dec        r5, r5
304=>x"BE6C",   -- 1011111001101100  brine      r5, mult_16_16.loop
305=>x"E383",   -- 1110001110000011  ba -, r6

306=>x"2449",   -- 0010010001001001  xor        r1, r1, r1
307=>x"C084",   -- 1100000010000100  li r4, 16
308=>x"0800",   -- 0000100000000000  add        r0, r0, r0
309=>x"0C49",   -- 0000110001001001  adc        r1, r1, r1
310=>x"0A8B",   -- 0000101010001011  sub        r3, r1, r2
311=>x"80DD",   -- 1000000011011101  brilt      r3, div_16_16.skip
312=>x"0A89",   -- 0000101010001001  sub        r1, r1, r2
313=>x"0400",   -- 0000010000000000  inc        r0, r0
314=>x"0624",   -- 0000011000100100  dec        r4, r4
315=>x"BE64",   -- 1011111001100100  brine      r4, div_16_16.loop
316=>x"E383",   -- 1110001110000011  ba -, r6

317=>x"2400",   -- 0010010000000000  xor        r0, r0, r0
318=>x"2449",   -- 0010010001001001  xor        r1, r1, r1
319=>x"8250",   -- 1000001001010000  brieq      r2, fact_16.end
320=>x"0409",   -- 0000010000001001  inc        r1, r1
321=>x"1008",   -- 0001000000001000  mova       r0, r1
322=>x"FAF0",   -- 1111101011110000  bail       -, r6, mult_16_16
323=>x"0126",   -- 0000000100100110  
324=>x"8104",   -- 1000000100000100  brine      r0, fact_16.overflow
325=>x"0126",   -- 0000000100100110  
326=>x"0612",   -- 0000011000010010  dec        r2, r2
327=>x"BE94",   -- 1011111010010100  brine      r2, fact_16.loop
328=>x"E383",   -- 1110001110000011  ba -, r6

329=>x"460C",   -- 0100011000001100  shl r4, r1, 3
330=>x"4209",   -- 0100001000001001  shl        r1, r1, 1
331=>x"0864",   -- 0000100001100100  add        r4, r4, r1
332=>x"0824",   -- 0000100000100100  add        r4, r4, r0
333=>x"D011",   -- 1101000000010001  lw r1, r2
334=>x"D221",   -- 1101001000100001  sw r1, r4
335=>x"0412",   -- 0000010000010010  inc        r2, r2
336=>x"0424",   -- 0000010000100100  inc        r4, r4
337=>x"061B",   -- 0000011000011011  dec        r3, r3
338=>x"BEDC",   -- 1011111011011100  brine      r3, put_sprite_16_aligned.loop
339=>x"E383",   -- 1110001110000011  ba -, r6

340=>x"460C",   -- 0100011000001100  shl r4, r1, 3
341=>x"4209",   -- 0100001000001001  shl        r1, r1, 1
342=>x"0864",   -- 0000100001100100  add        r4, r4, r1
343=>x"4001",   -- 0100000000000001  shl        r1, r0, 0
344=>x"0E00",   -- 0000111000000000  sbc        r0, r0, r0
345=>x"0864",   -- 0000100001100100  add        r4, r4, r1
346=>x"C0A5",   -- 1100000010100101  li r5, 20
347=>x"83C4",   -- 1000001111000100  brine      r0, put_sprite_8_aligned.loop1
348=>x"D010",   -- 1101000000010000  lw r0, r2
349=>x"D021",   -- 1101000000100001  lw r1, r4
350=>x"1A41",   -- 0001101001000001  mixhl      r1, r0, r1
351=>x"D221",   -- 1101001000100001  sw r1, r4
352=>x"061B",   -- 0000011000011011  dec        r3, r3
353=>x"8218",   -- 1000001000011000  brieq      r3, put_sprite_8_aligned.end
354=>x"0964",   -- 0000100101100100  add        r4, r4, r5
355=>x"D021",   -- 1101000000100001  lw r1, r4
356=>x"1E41",   -- 0001111001000001  mixll      r1, r0, r1
357=>x"D221",   -- 1101001000100001  sw r1, r4
358=>x"0412",   -- 0000010000010010  inc        r2, r2
359=>x"061B",   -- 0000011000011011  dec        r3, r3
360=>x"BD1C",   -- 1011110100011100  brine      r3, put_sprite_8_aligned.loop0
361=>x"E383",   -- 1110001110000011  ba -, r6
362=>x"D010",   -- 1101000000010000  lw r0, r2
363=>x"D021",   -- 1101000000100001  lw r1, r4
364=>x"1809",   -- 0001100000001001  mixhh      r1, r1, r0
365=>x"D221",   -- 1101001000100001  sw r1, r4
366=>x"061B",   -- 0000011000011011  dec        r3, r3
367=>x"BE98",   -- 1011111010011000  brieq      r3, put_sprite_8_aligned.end
368=>x"0964",   -- 0000100101100100  add        r4, r4, r5
369=>x"D021",   -- 1101000000100001  lw r1, r4
370=>x"1A09",   -- 0001101000001001  mixhl      r1, r1, r0
371=>x"D221",   -- 1101001000100001  sw r1, r4
372=>x"0412",   -- 0000010000010010  inc        r2, r2
373=>x"061B",   -- 0000011000011011  dec        r3, r3
374=>x"BD1C",   -- 1011110100011100  brine      r3, put_sprite_8_aligned.loop1
375=>x"E383",   -- 1110001110000011  ba -, r6

--     0=>X"D400", -- IN R0
--     1=>X"D600", -- OUT R0
--     2=>X"8043", -- bri r0, 1
--     3=>X"D400", -- IN R0
--     4=>X"D600", -- OUT R0
--     5=>X"FFFF", -- RESET
    others => x"0000"
    );
begin
  process(CLK)
  begin
    if (CLK'event AND CLK='1') then
      D <= m(to_integer(unsigned(AD)));
    end if;
  end process;
end Behavioral;
