----------------------------------------------------------------------------------
--
-- File retrieved, on 07/02/2010, from :
-- http://sebastien-viardot.imag.fr/Enseignements/Archi1A2s/sources/ROMPROG.vhd
--
-- Slightly altered to get rid of vendor-specific packages and adjust formatting
-- Now auto-filled by asrom script
--
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROMPROG is
  Port ( AD : in  STD_LOGIC_VECTOR (12 downto 0);
         D : out  STD_LOGIC_VECTOR (15 downto 0);
         CLK : in STD_LOGIC);
end ROMPROG;

architecture Behavioral of ROMPROG is
  constant low_address: natural := 0;
  constant high_address: natural := 8192;
  subtype octet is std_logic_vector( 15 downto 0 );
  type zone_memoire is
    array (natural range low_address to high_address-1) of octet;
  constant m: zone_memoire:= (
    0=>x"FFF7",	-- 1111111111110111  liw	r7, IRQ_mask
    1=>x"2000",	-- 0010000000000000  
    2=>x"F8C0",	-- 1111100011000000  bai	-, os_init
    3=>x"0100",	-- 0000000100000000  
   16=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_ack
   17=>x"2002",	-- 0010000000000010  
   18=>x"D001",	-- 1101000000000001  lw	r1, r0
   19=>x"F54A",	-- 1111010101001010  bspl	r2, r1, 5
   20=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_error
   21=>x"00A0",	-- 0000000010100000  
   22=>x"F4CA",	-- 1111010011001010  bspl	r2, r1, 3
   23=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_kbd
   24=>x"0090",	-- 0000000010010000  
   25=>x"F40A",	-- 1111010000001010  bspl	r2, r1, 0
   26=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_tmr
   27=>x"0080",	-- 0000000010000000  
   28=>x"CFF9",	-- 1100111111111001  li	r1, -1
   29=>x"D201",	-- 1101001000000001  sw	r1, r0
   30=>x"FFFE",	-- 1111111111111110  reti
  128=>x"2624",	-- 0010011000100100  not r4, r4
  129=>x"D700",	-- 1101011100000000  out	r4
  130=>x"E383",	-- 1110001110000011  ba	-, r6
  144=>x"E383",	-- 1110001110000011  ba	-, r6
  160=>x"2524",	-- 0010010100100100  xor	r4, r4, r4
  161=>x"D700",	-- 1101011100000000  out	r4
  162=>x"E383",	-- 1110001110000011  ba	-, r6
  256=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_mask
  257=>x"2000",	-- 0010000000000000  
  258=>x"C0C9",	-- 1100000011001001  li	r1, 0x19
  259=>x"D201",	-- 1101001000000001  sw	r1, r0
  260=>x"0400",	-- 0000010000000000  inc	r0, r0
  261=>x"CFF9",	-- 1100111111111001  li	r1, -1
  262=>x"D201",	-- 1101001000000001  sw	r1, r0
  263=>x"C03A",	-- 1100000000111010  li	r2, 7
  264=>x"0880",	-- 0000100010000000  add	r0, r0, r2
  265=>x"C0EA",	-- 1100000011101010  li	r2, 0x1D
  266=>x"D202",	-- 1101001000000010  sw	r2, r0
  267=>x"0400",	-- 0000010000000000  inc	r0, r0
  268=>x"C07A",	-- 1100000001111010  li	r2, 15
  269=>x"D202",	-- 1101001000000010  sw	r2, r0
  270=>x"FFF0",	-- 1111111111110000  liw	r0, 0x8421
  271=>x"8421",	-- 1000010000100001  
  272=>x"FFF1",	-- 1111111111110001  liw	r1, 0x1234
  273=>x"1234",	-- 0001001000110100  
  274=>x"D640",	-- 1101011001000000  out	r1
  275=>x"E408",	-- 1110010000001000  exw	r0, r1
  276=>x"E408",	-- 1110010000001000  exw	r0, r1
  277=>x"1842",	-- 0001100001000010  mixhh	r2, r0, r1
  278=>x"1A43",	-- 0001101001000011  mixhl	r3, r0, r1
  279=>x"1C44",	-- 0001110001000100  mixlh	r4, r0, r1
  280=>x"1E45",	-- 0001111001000101  mixll	r5, r0, r1
  281=>x"C01E",	-- 1100000000011110  li	r6, 3
  282=>x"3985",	-- 0011100110000101  rrr	r5, r0, r6
  283=>x"3B8D",	-- 0011101110001101  rrl	r5, r1, r6
  284=>x"3D95",	-- 0011110110010101  rsr	r5, r2, r6
  285=>x"3F9D",	-- 0011111110011101  rsl	r5, r3, r6
  286=>x"FC0E",	-- 1111110000001110  mul	r6, r1, r0
  287=>x"C028",	-- 1100000000101000  li	r0, 5
  288=>x"C151",	-- 1100000101010001  li	r1, 42
  289=>x"FFF2",	-- 1111111111110010  liw	r2, font_map + 4 * 0x23
  290=>x"134C",	-- 0001001101001100  
  291=>x"C043",	-- 1100000001000011  li	r3, 8
  292=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  293=>x"01E5",	-- 0000000111100101  
  294=>x"C000",	-- 1100000000000000  li	r0, 0
  295=>x"C0A1",	-- 1100000010100001  li	r1, 20
  296=>x"FFF2",	-- 1111111111110010  liw	r2, hello_str
  297=>x"16C0",	-- 0001011011000000  
  298=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  299=>x"01A5",	-- 0000000110100101  
  300=>x"2400",	-- 0010010000000000  xor	r0, r0, r0
  301=>x"C0A1",	-- 1100000010100001  li	r1, 20
  302=>x"FFF2",	-- 1111111111110010  liw	r2, 0x2020
  303=>x"2020",	-- 0010000000100000  
  304=>x"D202",	-- 1101001000000010  sw	r2, r0
  305=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  306=>x"FFF2",	-- 1111111111110010  liw	r2, 0x7070
  307=>x"7070",	-- 0111000001110000  
  308=>x"D202",	-- 1101001000000010  sw	r2, r0
  309=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  310=>x"FFF2",	-- 1111111111110010  liw	r2, 0xF8F8
  311=>x"F8F8",	-- 1111100011111000  
  312=>x"D202",	-- 1101001000000010  sw	r2, r0
  313=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  314=>x"FFF2",	-- 1111111111110010  liw	r2, 0xF8F8
  315=>x"F8F8",	-- 1111100011111000  
  316=>x"D202",	-- 1101001000000010  sw	r2, r0
  317=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  318=>x"FFF2",	-- 1111111111110010  liw	r2, 0xF870
  319=>x"F870",	-- 1111100001110000  
  320=>x"D202",	-- 1101001000000010  sw	r2, r0
  321=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  322=>x"FFF2",	-- 1111111111110010  liw	r2, 0x7020
  323=>x"7020",	-- 0111000000100000  
  324=>x"D202",	-- 1101001000000010  sw	r2, r0
  325=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  326=>x"FFF2",	-- 1111111111110010  liw	r2, 0x2070
  327=>x"2070",	-- 0010000001110000  
  328=>x"D202",	-- 1101001000000010  sw	r2, r0
  329=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  330=>x"FFF2",	-- 1111111111110010  liw	r2, 0x0000
  332=>x"D202",	-- 1101001000000010  sw	r2, r0
  333=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  334=>x"C000",	-- 1100000000000000  li	r0, 0
  335=>x"C0F1",	-- 1100000011110001  li	r1, 30
  336=>x"FFF2",	-- 1111111111110010  liw	r2, font_map
  337=>x"12C0",	-- 0001001011000000  
  338=>x"FFF3",	-- 1111111111110011  liw	r3, PS2_stat
  339=>x"2006",	-- 0010000000000110  
  340=>x"D01B",	-- 1101000000011011  lw	r3, r3
  341=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  342=>x"87E4",	-- 1000011111100100  brine	r4, event_not_kbd
  343=>x"063F",	-- 0000011000111111  dec	r7, r7
  344=>x"D23A",	-- 1101001000111010  sw	r2, r7
  345=>x"063F",	-- 0000011000111111  dec	r7, r7
  346=>x"D238",	-- 1101001000111000  sw	r0, r7
  347=>x"063F",	-- 0000011000111111  dec	r7, r7
  348=>x"D239",	-- 1101001000111001  sw	r1, r7
  349=>x"FFF3",	-- 1111111111110011  liw	r3, PS2_rx
  350=>x"2004",	-- 0010000000000100  
  351=>x"D01B",	-- 1101000000011011  lw	r3, r3
  352=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  353=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  354=>x"C043",	-- 1100000001000011  li	r3, 8
  355=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  356=>x"01E5",	-- 0000000111100101  
  357=>x"D039",	-- 1101000000111001  lw	r1, r7
  358=>x"043F",	-- 0000010000111111  inc	r7, r7
  359=>x"D038",	-- 1101000000111000  lw	r0, r7
  360=>x"043F",	-- 0000010000111111  inc	r7, r7
  361=>x"0400",	-- 0000010000000000  inc	r0, r0
  362=>x"C142",	-- 1100000101000010  li	r2, 40
  363=>x"0A82",	-- 0000101010000010  sub	r2, r0, r2
  364=>x"81D5",	-- 1000000111010101  brilt	r2, event_kbd_end
  365=>x"C042",	-- 1100000001000010  li	r2, 8
  366=>x"0889",	-- 0000100010001001  add	r1, r1, r2
  367=>x"C74A",	-- 1100011101001010  li	r2, 233
  368=>x"0A8A",	-- 0000101010001010  sub	r2, r1, r2
  369=>x"8095",	-- 1000000010010101  brilt	r2, event_kbd_end
  370=>x"C0F1",	-- 1100000011110001  li	r1, 30
  371=>x"D03A",	-- 1101000000111010  lw	r2, r7
  372=>x"043F",	-- 0000010000111111  inc	r7, r7
  373=>x"B743",	-- 1011011101000011  bri	-, event_loop
  374=>x"C750",	-- 1100011101010000  li	r0, 234
  375=>x"C1C2",	-- 1100000111000010  li	r2, 56
  376=>x"FAC6",	-- 1111101011000110  bail	-, r6, div_16_16
  377=>x"018E",	-- 0000000110001110  
  378=>x"C448",	-- 1100010001001000  li	r0, 137
  379=>x"C472",	-- 1100010001110010  li	r2, 142
  380=>x"FAC6",	-- 1111101011000110  bail	-, r6, mult_16_16
  381=>x"0182",	-- 0000000110000010  
  382=>x"C03A",	-- 1100000000111010  li r2, 7
  383=>x"FAC6",	-- 1111101011000110  bail	-, r6, fact_16
  384=>x"0199",	-- 0000000110011001  
  385=>x"FFFF",	-- 1111111111111111  reset
  386=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  387=>x"2524",	-- 0010010100100100  xor	r4, r4, r4
  388=>x"C085",	-- 1100000010000101  li	r5, 16
  389=>x"0849",	-- 0000100001001001  add	r1, r1, r1
  390=>x"0C00",	-- 0000110000000000  adc	r0, r0, r0
  391=>x"0EDB",	-- 0000111011011011  sbc	r3, r3, r3
  392=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  393=>x"08C9",	-- 0000100011001001  add	r1, r1, r3
  394=>x"0D00",	-- 0000110100000000  adc	r0, r0, r4
  395=>x"062D",	-- 0000011000101101  dec	r5, r5
  396=>x"BE6C",	-- 1011111001101100  brine	r5, mult_16_16.loop
  397=>x"E383",	-- 1110001110000011  ba	-, r6
  398=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  399=>x"C084",	-- 1100000010000100  li	r4, 16
  400=>x"0800",	-- 0000100000000000  add	r0, r0, r0
  401=>x"0C49",	-- 0000110001001001  adc	r1, r1, r1
  402=>x"0A8B",	-- 0000101010001011  sub	r3, r1, r2
  403=>x"80DD",	-- 1000000011011101  brilt	r3, div_16_16.skip
  404=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  405=>x"0400",	-- 0000010000000000  inc	r0, r0
  406=>x"0624",	-- 0000011000100100  dec	r4, r4
  407=>x"BE64",	-- 1011111001100100  brine	r4, div_16_16.loop
  408=>x"E383",	-- 1110001110000011  ba	-, r6
  409=>x"2400",	-- 0010010000000000  xor	r0, r0, r0
  410=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  411=>x"8250",	-- 1000001001010000  brieq	r2, fact_16.end
  412=>x"0409",	-- 0000010000001001  inc	r1, r1
  413=>x"1008",	-- 0001000000001000  mova	r0, r1
  414=>x"FAC6",	-- 1111101011000110  bail	-, r6, mult_16_16
  415=>x"0182",	-- 0000000110000010  
  416=>x"8104",	-- 1000000100000100  brine	r0, fact_16.overflow
  417=>x"0182",	-- 0000000110000010  
  418=>x"0612",	-- 0000011000010010  dec	r2, r2
  419=>x"BE94",	-- 1011111010010100  brine	r2, fact_16.loop
  420=>x"E383",	-- 1110001110000011  ba	-, r6
  421=>x"063F",	-- 0000011000111111  dec	r7, r7
  422=>x"D23E",	-- 1101001000111110  sw	r6, r7
  423=>x"D013",	-- 1101000000010011  lw	r3, r2
  424=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  425=>x"8B98",	-- 1000101110011000  brieq	r3, puts.end
  426=>x"063F",	-- 0000011000111111  dec	r7, r7
  427=>x"D238",	-- 1101001000111000  sw	r0, r7
  428=>x"063F",	-- 0000011000111111  dec	r7, r7
  429=>x"D239",	-- 1101001000111001  sw	r1, r7
  430=>x"063F",	-- 0000011000111111  dec	r7, r7
  431=>x"D23A",	-- 1101001000111010  sw	r2, r7
  432=>x"FFF4",	-- 1111111111110100  liw	r4, font_map
  433=>x"12C0",	-- 0001001011000000  
  434=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  435=>x"091A",	-- 0000100100011010  add	r2, r3, r4
  436=>x"C043",	-- 1100000001000011  li	r3, 8
  437=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  438=>x"01E5",	-- 0000000111100101  
  439=>x"D03A",	-- 1101000000111010  lw	r2, r7
  440=>x"043F",	-- 0000010000111111  inc	r7, r7
  441=>x"D039",	-- 1101000000111001  lw	r1, r7
  442=>x"043F",	-- 0000010000111111  inc	r7, r7
  443=>x"D038",	-- 1101000000111000  lw	r0, r7
  444=>x"043F",	-- 0000010000111111  inc	r7, r7
  445=>x"0400",	-- 0000010000000000  inc	r0, r0
  446=>x"D013",	-- 1101000000010011  lw	r3, r2
  447=>x"4E1B",	-- 0100111000011011  shl	r3, r3, 7
  448=>x"6A1B",	-- 0110101000011011  shr	r3, r3, 5
  449=>x"8598",	-- 1000010110011000  brieq	r3, puts.end
  450=>x"063F",	-- 0000011000111111  dec	r7, r7
  451=>x"D238",	-- 1101001000111000  sw	r0, r7
  452=>x"063F",	-- 0000011000111111  dec	r7, r7
  453=>x"D239",	-- 1101001000111001  sw	r1, r7
  454=>x"063F",	-- 0000011000111111  dec	r7, r7
  455=>x"D23A",	-- 1101001000111010  sw	r2, r7
  456=>x"FFF4",	-- 1111111111110100  liw	r4, font_map
  457=>x"12C0",	-- 0001001011000000  
  458=>x"091A",	-- 0000100100011010  add	r2, r3, r4
  459=>x"C043",	-- 1100000001000011  li	r3, 8
  460=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  461=>x"01E5",	-- 0000000111100101  
  462=>x"D03A",	-- 1101000000111010  lw	r2, r7
  463=>x"043F",	-- 0000010000111111  inc	r7, r7
  464=>x"D039",	-- 1101000000111001  lw	r1, r7
  465=>x"043F",	-- 0000010000111111  inc	r7, r7
  466=>x"D038",	-- 1101000000111000  lw	r0, r7
  467=>x"043F",	-- 0000010000111111  inc	r7, r7
  468=>x"0400",	-- 0000010000000000  inc	r0, r0
  469=>x"0412",	-- 0000010000010010  inc	r2, r2
  470=>x"B443",	-- 1011010001000011  bri	-, puts.loop
  471=>x"D03E",	-- 1101000000111110  lw	r6, r7
  472=>x"043F",	-- 0000010000111111  inc	r7, r7
  473=>x"E383",	-- 1110001110000011  ba	-, r6
  474=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  475=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  476=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  477=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  478=>x"D011",	-- 1101000000010001  lw	r1, r2
  479=>x"D221",	-- 1101001000100001  sw	r1, r4
  480=>x"0412",	-- 0000010000010010  inc	r2, r2
  481=>x"0424",	-- 0000010000100100  inc	r4, r4
  482=>x"061B",	-- 0000011000011011  dec	r3, r3
  483=>x"BEDC",	-- 1011111011011100  brine	r3, put_sprite_16_aligned.loop
  484=>x"E383",	-- 1110001110000011  ba	-, r6
  485=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  486=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  487=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  488=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  489=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  490=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  491=>x"C0A5",	-- 1100000010100101  li	r5, 20
  492=>x"8404",	-- 1000010000000100  brine	r0, put_sprite_8_aligned.loop1
  493=>x"D010",	-- 1101000000010000  lw	r0, r2
  494=>x"D021",	-- 1101000000100001  lw	r1, r4
  495=>x"1A41",	-- 0001101001000001  mixhl	r1, r0, r1
  496=>x"D221",	-- 1101001000100001  sw	r1, r4
  497=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  498=>x"061B",	-- 0000011000011011  dec	r3, r3
  499=>x"E398",	-- 1110001110011000  baeq	r3, r6
  500=>x"D021",	-- 1101000000100001  lw	r1, r4
  501=>x"1E41",	-- 0001111001000001  mixll	r1, r0, r1
  502=>x"D221",	-- 1101001000100001  sw	r1, r4
  503=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  504=>x"0412",	-- 0000010000010010  inc	r2, r2
  505=>x"061B",	-- 0000011000011011  dec	r3, r3
  506=>x"E398",	-- 1110001110011000  baeq	r3, r6
  507=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop0
  508=>x"D010",	-- 1101000000010000  lw	r0, r2
  509=>x"D021",	-- 1101000000100001  lw	r1, r4
  510=>x"1809",	-- 0001100000001001  mixhh	r1, r1, r0
  511=>x"D221",	-- 1101001000100001  sw	r1, r4
  512=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  513=>x"061B",	-- 0000011000011011  dec	r3, r3
  514=>x"E398",	-- 1110001110011000  baeq	r3, r6
  515=>x"D021",	-- 1101000000100001  lw	r1, r4
  516=>x"1A09",	-- 0001101000001001  mixhl	r1, r1, r0
  517=>x"D221",	-- 1101001000100001  sw	r1, r4
  518=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  519=>x"0412",	-- 0000010000010010  inc	r2, r2
  520=>x"061B",	-- 0000011000011011  dec	r3, r3
  521=>x"E398",	-- 1110001110011000  baeq	r3, r6
  522=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop1
    others => x"0000"
    );
begin
  process(CLK)
  begin
    if (CLK'event AND CLK='1') then
      D <= m(to_integer(unsigned(AD)));
    end if;
  end process;
end Behavioral;
