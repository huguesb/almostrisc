----------------------------------------------------------------------------------
--
-- File retrieved, on 07/02/2010, from :
-- http://sebastien-viardot.imag.fr/Enseignements/Archi1A2s/sources/ROMPROG.vhd
--
-- Slightly altered to get rid of vendor-specific packages and adjust formatting
-- Now auto-filled by asrom script
--
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROMPROG is
  Port ( AD : in  STD_LOGIC_VECTOR (12 downto 0);
         D : out  STD_LOGIC_VECTOR (15 downto 0);
         CLK : in STD_LOGIC);
end ROMPROG;

architecture Behavioral of ROMPROG is
  constant low_address: natural := 0;
  constant high_address: natural := 8192;
  subtype octet is std_logic_vector( 15 downto 0 );
  type zone_memoire is
    array (natural range low_address to high_address-1) of octet;
  constant m: zone_memoire:= (
    0=>x"FFF7",	-- 1111111111110111  liw	r7, IRQ_mask
    1=>x"2000",	-- 0010000000000000  
    2=>x"F8C0",	-- 1111100011000000  bai	-, os_init
    3=>x"0100",	-- 0000000100000000  
   16=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_ack
   17=>x"2002",	-- 0010000000000010  
   18=>x"D001",	-- 1101000000000001  lw	r1, r0
   19=>x"F54A",	-- 1111010101001010  bspl	r2, r1, 5
   20=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_error
   21=>x"0050",	-- 0000000001010000  
   22=>x"F4CA",	-- 1111010011001010  bspl	r2, r1, 3
   23=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_kbd
   24=>x"0060",	-- 0000000001100000  
   25=>x"F40A",	-- 1111010000001010  bspl	r2, r1, 0
   26=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_tmr
   27=>x"0040",	-- 0000000001000000  
   28=>x"D201",	-- 1101001000000001  sw	r1, r0
   29=>x"FFFE",	-- 1111111111111110  reti
   64=>x"263F",	-- 0010011000111111  not r7, r7
   65=>x"D7C0",	-- 1101011111000000  out	r7
   66=>x"E383",	-- 1110001110000011  ba	-, r6
   80=>x"25FF",	-- 0010010111111111  xor	r7, r7, r7
   81=>x"D7C0",	-- 1101011111000000  out	r7
   82=>x"E383",	-- 1110001110000011  ba	-, r6
   96=>x"FFF2",	-- 1111111111110010  liw	r2, PS2_rx
   97=>x"2004",	-- 0010000000000100  
   98=>x"D012",	-- 1101000000010010  lw	r2, r2
   99=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map + 8
  100=>x"1808",	-- 0001100000001000  
  101=>x"D01B",	-- 1101000000011011  lw	r3, r3
  102=>x"1EBF",	-- 0001111010111111  mixll	r7, r7, r2
  103=>x"C784",	-- 1100011110000100  li	r4, 0xF0
  104=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  105=>x"8B20",	-- 1000101100100000  brieq	r4, int_kbd.release
  106=>x"C704",	-- 1100011100000100  li	r4, 0xE0
  107=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  108=>x"88E0",	-- 1000100011100000  brieq	r4, int_kbd.extended
  109=>x"FFF5",	-- 1111111111110101  liw	r5, 0x16C0 - 1
  110=>x"16BF",	-- 0001011010111111  
  111=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  112=>x"80E0",	-- 1000000011100000  brieq	r4, $+3
  113=>x"FFF5",	-- 1111111111110101  liw	r5, 0x16CA - 1
  114=>x"16C9",	-- 0001011011001001  
  115=>x"042D",	-- 0000010000101101  inc	r5, r5
  116=>x"D02C",	-- 1101000000101100  lw	r4, r5
  117=>x"8560",	-- 1000010101100000  brieq	r4, scan_code_mismatch
  118=>x"6E24",	-- 0110111000100100  shr	r4, r4, 7
  119=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  120=>x"BEE4",	-- 1011111011100100  brine	r4, scan_code_loop
  121=>x"D02A",	-- 1101000000101010  lw	r2, r5
  122=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  123=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  124=>x"741B",	-- 0111010000011011  shr	r3, r3, 10
  125=>x"C00D",	-- 1100000000001101  li	r5, 1
  126=>x"0612",	-- 0000011000010010  dec	r2, r2
  127=>x"3AAA",	-- 0011101010101010  rrl	r2, r5, r2
  128=>x"FFF5",	-- 1111111111110101  liw	r5, key_press_map
  129=>x"1800",	-- 0001100000000000  
  130=>x"08ED",	-- 0000100011101101  add	r5, r5, r3
  131=>x"D02B",	-- 1101000000101011  lw	r3, r5
  132=>x"80E4",	-- 1000000011100100  brine	r4, scan_code_release
  133=>x"229B",	-- 0010001010011011  or	r3, r3, r2
  134=>x"80C3",	-- 1000000011000011  bri	-, scan_code_notify
  135=>x"2612",	-- 0010011000010010  not	r2, r2
  136=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  137=>x"D22B",	-- 1101001000101011  sw	r3, r5
  138=>x"C003",	-- 1100000000000011  li	r3, 0
  139=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  140=>x"1808",	-- 0001100000001000  
  141=>x"D223",	-- 1101001000100011  sw	r3, r4
  142=>x"E383",	-- 1110001110000011  ba	-, r6
  143=>x"C014",	-- 1100000000010100  li	r4, 2
  144=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  145=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  146=>x"1808",	-- 0001100000001000  
  147=>x"D223",	-- 1101001000100011  sw	r3, r4
  148=>x"E383",	-- 1110001110000011  ba	-, r6
  149=>x"C00C",	-- 1100000000001100  li	r4, 1
  150=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  151=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  152=>x"1808",	-- 0001100000001000  
  153=>x"D223",	-- 1101001000100011  sw	r3, r4
  154=>x"E383",	-- 1110001110000011  ba	-, r6
  256=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_mask
  257=>x"2000",	-- 0010000000000000  
  258=>x"C0C9",	-- 1100000011001001  li	r1, 0x19
  259=>x"D201",	-- 1101001000000001  sw	r1, r0
  260=>x"0400",	-- 0000010000000000  inc	r0, r0
  261=>x"CFF9",	-- 1100111111111001  li	r1, -1
  262=>x"D201",	-- 1101001000000001  sw	r1, r0
  263=>x"C03A",	-- 1100000000111010  li	r2, 7
  264=>x"0880",	-- 0000100010000000  add	r0, r0, r2
  265=>x"C0EA",	-- 1100000011101010  li	r2, 0x1D
  266=>x"D202",	-- 1101001000000010  sw	r2, r0
  267=>x"0400",	-- 0000010000000000  inc	r0, r0
  268=>x"C07A",	-- 1100000001111010  li	r2, 15
  269=>x"D202",	-- 1101001000000010  sw	r2, r0
  270=>x"FFF0",	-- 1111111111110000  liw	r0, key_press_map
  271=>x"1800",	-- 0001100000000000  
  272=>x"C001",	-- 1100000000000001  li	r1, 0
  273=>x"C042",	-- 1100000001000010  li	r2, 8
  274=>x"D201",	-- 1101001000000001  sw	r1, r0
  275=>x"0400",	-- 0000010000000000  inc	r0, r0
  276=>x"0612",	-- 0000011000010010  dec	r2, r2
  277=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  278=>x"C0F3",	-- 1100000011110011  li	r3, 30
  279=>x"CFFA",	-- 1100111111111010  li	r2, -1
  280=>x"D21A",	-- 1101001000011010  sw	r2, r3
  281=>x"8083",	-- 1000000010000011  bri	-, PaperGameStart
  282=>x"8003",	-- 1000000000000011  bri	-, PaperMenuLoop
  283=>x"C000",	-- 1100000000000000  li	r0, 0
  284=>x"FFF1",	-- 1111111111110001  liw	r1, 0x0801
  285=>x"0801",	-- 0000100000000001  
  286=>x"063F",	-- 0000011000111111  dec	r7, r7
  287=>x"D238",	-- 1101001000111000  sw	r0, r7
  288=>x"063F",	-- 0000011000111111  dec	r7, r7
  289=>x"D239",	-- 1101001000111001  sw	r1, r7
  290=>x"063F",	-- 0000011000111111  dec	r7, r7
  291=>x"D23A",	-- 1101001000111010  sw	r2, r7
  292=>x"C000",	-- 1100000000000000  li	r0, 0
  293=>x"CFF9",	-- 1100111111111001  li	r1, -1
  294=>x"C0A2",	-- 1100000010100010  li	r2, 20
  295=>x"D201",	-- 1101001000000001  sw	r1, r0
  296=>x"0400",	-- 0000010000000000  inc	r0, r0
  297=>x"0612",	-- 0000011000010010  dec	r2, r2
  298=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  299=>x"C001",	-- 1100000000000001  li	r1, 0
  300=>x"FFF2",	-- 1111111111110010  liw	r2, 18*20
  301=>x"0168",	-- 0000000101101000  
  302=>x"D201",	-- 1101001000000001  sw	r1, r0
  303=>x"0400",	-- 0000010000000000  inc	r0, r0
  304=>x"0612",	-- 0000011000010010  dec	r2, r2
  305=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  306=>x"CFF9",	-- 1100111111111001  li	r1, -1
  307=>x"C0A2",	-- 1100000010100010  li	r2, 20
  308=>x"D201",	-- 1101001000000001  sw	r1, r0
  309=>x"0400",	-- 0000010000000000  inc	r0, r0
  310=>x"0612",	-- 0000011000010010  dec	r2, r2
  311=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  312=>x"C020",	-- 1100000000100000  li	r0, 4
  313=>x"C029",	-- 1100000000101001  li	r1, 5
  314=>x"FFF2",	-- 1111111111110010  liw	r2, paper_title
  315=>x"1730",	-- 0001011100110000  
  316=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  317=>x"01F8",	-- 0000000111111000  
  318=>x"C790",	-- 1100011110010000  li	r0, 242
  319=>x"C009",	-- 1100000000001001  li	r1, 1
  320=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud
  321=>x"1720",	-- 0001011100100000  
  322=>x"C043",	-- 1100000001000011  li	r3, 8
  323=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  324=>x"0283",	-- 0000001010000011  
  325=>x"C118",	-- 1100000100011000  li	r0, 35
  326=>x"C009",	-- 1100000000001001  li	r1, 1
  327=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  328=>x"1736",	-- 0001011100110110  
  329=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  330=>x"01F8",	-- 0000000111111000  
  331=>x"C790",	-- 1100011110010000  li	r0, 242
  332=>x"C051",	-- 1100000001010001  li	r1, 10
  333=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud + 4
  334=>x"1724",	-- 0001011100100100  
  335=>x"C043",	-- 1100000001000011  li	r3, 8
  336=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  337=>x"0283",	-- 0000001010000011  
  338=>x"C118",	-- 1100000100011000  li	r0, 35
  339=>x"C051",	-- 1100000001010001  li	r1, 10
  340=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  341=>x"1736",	-- 0001011100110110  
  342=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  343=>x"01F8",	-- 0000000111111000  
  344=>x"D03A",	-- 1101000000111010  lw	r2, r7
  345=>x"043F",	-- 0000010000111111  inc	r7, r7
  346=>x"D039",	-- 1101000000111001  lw	r1, r7
  347=>x"043F",	-- 0000010000111111  inc	r7, r7
  348=>x"D038",	-- 1101000000111000  lw	r0, r7
  349=>x"043F",	-- 0000010000111111  inc	r7, r7
  350=>x"063F",	-- 0000011000111111  dec	r7, r7
  351=>x"D238",	-- 1101001000111000  sw	r0, r7
  352=>x"063F",	-- 0000011000111111  dec	r7, r7
  353=>x"D239",	-- 1101001000111001  sw	r1, r7
  354=>x"063F",	-- 0000011000111111  dec	r7, r7
  355=>x"D23A",	-- 1101001000111010  sw	r2, r7
  356=>x"C4C0",	-- 1100010011000000  li	r0, 152
  357=>x"C161",	-- 1100000101100001  li	r1, 44
  358=>x"FFF2",	-- 1111111111110010  liw	r2, paper_sprites
  359=>x"16D0",	-- 0001011011010000  
  360=>x"C083",	-- 1100000010000011  li	r3, 16
  361=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_16
  362=>x"0233",	-- 0000001000110011  
  363=>x"D03A",	-- 1101000000111010  lw	r2, r7
  364=>x"043F",	-- 0000010000111111  inc	r7, r7
  365=>x"D039",	-- 1101000000111001  lw	r1, r7
  366=>x"043F",	-- 0000010000111111  inc	r7, r7
  367=>x"D038",	-- 1101000000111000  lw	r0, r7
  368=>x"043F",	-- 0000010000111111  inc	r7, r7
  369=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  370=>x"1800",	-- 0001100000000000  
  371=>x"D01B",	-- 1101000000011011  lw	r3, r3
  372=>x"9518",	-- 1001010100011000  brieq	r3, event_not_kbd
  373=>x"F7DC",	-- 1111011111011100  bspl	r4, r3, 15
  374=>x"82A0",	-- 1000001010100000  brieq	r4, PaperGameQuit
  375=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  376=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveUp
  377=>x"F49C",	-- 1111010010011100  bspl	r4, r3, 2
  378=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveDOWN
  379=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  380=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveLEFT
  381=>x"F4DC",	-- 1111010011011100  bspl	r4, r3, 3
  382=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveRIGHT
  383=>x"BC83",	-- 1011110010000011  bri	-, PaperGameLoop
  384=>x"FFFF",	-- 1111111111111111  reset
  385=>x"C040",	-- 1100000001000000  li	r0, 8
  386=>x"C041",	-- 1100000001000001  li	r1, 8
  387=>x"063F",	-- 0000011000111111  dec	r7, r7
  388=>x"D239",	-- 1101001000111001  sw	r1, r7
  389=>x"063F",	-- 0000011000111111  dec	r7, r7
  390=>x"D238",	-- 1101001000111000  sw	r0, r7
  391=>x"FFF2",	-- 1111111111110010  liw	r2, font_map + 4 * 0x23
  392=>x"134C",	-- 0001001101001100  
  393=>x"C043",	-- 1100000001000011  li	r3, 8
  394=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  395=>x"0283",	-- 0000001010000011  
  396=>x"D038",	-- 1101000000111000  lw	r0, r7
  397=>x"043F",	-- 0000010000111111  inc	r7, r7
  398=>x"D039",	-- 1101000000111001  lw	r1, r7
  399=>x"043F",	-- 0000010000111111  inc	r7, r7
  400=>x"C0A2",	-- 1100000010100010  li	r2, 20
  401=>x"C003",	-- 1100000000000011  li	r3, 0
  402=>x"061B",	-- 0000011000011011  dec	r3, r3
  403=>x"BFDC",	-- 1011111111011100  brine	r3, $-1
  404=>x"0612",	-- 0000011000010010  dec	r2, r2
  405=>x"BF14",	-- 1011111100010100  brine	r2, $-4
  406=>x"FFF2",	-- 1111111111110010  liw	r2, key_press_map
  407=>x"1800",	-- 0001100000000000  
  408=>x"D012",	-- 1101000000010010  lw	r2, r2
  409=>x"8BD0",	-- 1000101111010000  brieq	r2, event_not_kbd
  410=>x"063F",	-- 0000011000111111  dec	r7, r7
  411=>x"D23A",	-- 1101001000111010  sw	r2, r7
  412=>x"063F",	-- 0000011000111111  dec	r7, r7
  413=>x"D239",	-- 1101001000111001  sw	r1, r7
  414=>x"063F",	-- 0000011000111111  dec	r7, r7
  415=>x"D238",	-- 1101001000111000  sw	r0, r7
  416=>x"FFF2",	-- 1111111111110010  liw	r2, font_map
  417=>x"12C0",	-- 0001001011000000  
  418=>x"C043",	-- 1100000001000011  li	r3, 8
  419=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  420=>x"0283",	-- 0000001010000011  
  421=>x"D038",	-- 1101000000111000  lw	r0, r7
  422=>x"043F",	-- 0000010000111111  inc	r7, r7
  423=>x"D039",	-- 1101000000111001  lw	r1, r7
  424=>x"043F",	-- 0000010000111111  inc	r7, r7
  425=>x"D03A",	-- 1101000000111010  lw	r2, r7
  426=>x"043F",	-- 0000010000111111  inc	r7, r7
  427=>x"F413",	-- 1111010000010011  bspl	r3, r2, 0
  428=>x"81D8",	-- 1000000111011000  brieq	r3, event_kbd_no_up
  429=>x"C043",	-- 1100000001000011  li	r3, 8
  430=>x"0ACB",	-- 0000101011001011  sub	r3, r1, r3
  431=>x"809C",	-- 1000000010011100  brine	r3, event_kbd_no_clip_up
  432=>x"C781",	-- 1100011110000001  li	r1, 240
  433=>x"C043",	-- 1100000001000011  li	r3, 8
  434=>x"0AC9",	-- 0000101011001001  sub	r1, r1, r3
  435=>x"F453",	-- 1111010001010011  bspl	r3, r2, 1
  436=>x"8118",	-- 1000000100011000  brieq	r3, event_kbd_no_left
  437=>x"8084",	-- 1000000010000100  brine	r0, event_kbd_no_clip_left
  438=>x"C9C0",	-- 1100100111000000  li	r0, 39*8
  439=>x"0600",	-- 0000011000000000  dec	r0, r0
  440=>x"F493",	-- 1111010010010011  bspl	r3, r2, 2
  441=>x"81D8",	-- 1000000111011000  brieq	r3, event_kbd_no_down
  442=>x"C743",	-- 1100011101000011  li	r3, 232
  443=>x"0ACB",	-- 0000101011001011  sub	r3, r1, r3
  444=>x"809D",	-- 1000000010011101  brilt	r3, event_kbd_no_clip_down
  445=>x"C001",	-- 1100000000000001  li	r1, 0
  446=>x"C043",	-- 1100000001000011  li	r3, 8
  447=>x"08C9",	-- 0000100011001001  add	r1, r1, r3
  448=>x"F4D3",	-- 1111010011010011  bspl	r3, r2, 3
  449=>x"8198",	-- 1000000110011000  brieq	r3, event_kbd_no_right
  450=>x"C9C3",	-- 1100100111000011  li	r3, 39*8
  451=>x"0AC3",	-- 0000101011000011  sub	r3, r0, r3
  452=>x"809D",	-- 1000000010011101  brilt	r3, event_kbd_no_clip_right
  453=>x"CFF8",	-- 1100111111111000  li	r0, -1
  454=>x"0400",	-- 0000010000000000  inc	r0, r0
  455=>x"AF03",	-- 1010111100000011  bri	-, redraw
  456=>x"B383",	-- 1011001110000011  bri	-, event_loop
  457=>x"C750",	-- 1100011101010000  li	r0, 234
  458=>x"C1C2",	-- 1100000111000010  li	r2, 56
  459=>x"FAC6",	-- 1111101011000110  bail	-, r6, div_16_16
  460=>x"01E1",	-- 0000000111100001  
  461=>x"C448",	-- 1100010001001000  li	r0, 137
  462=>x"C472",	-- 1100010001110010  li	r2, 142
  463=>x"FAC6",	-- 1111101011000110  bail	-, r6, mult_16_16
  464=>x"01D5",	-- 0000000111010101  
  465=>x"C03A",	-- 1100000000111010  li r2, 7
  466=>x"FAC6",	-- 1111101011000110  bail	-, r6, fact_16
  467=>x"01EC",	-- 0000000111101100  
  468=>x"FFFF",	-- 1111111111111111  reset
  469=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  470=>x"2524",	-- 0010010100100100  xor	r4, r4, r4
  471=>x"C085",	-- 1100000010000101  li	r5, 16
  472=>x"0849",	-- 0000100001001001  add	r1, r1, r1
  473=>x"0C00",	-- 0000110000000000  adc	r0, r0, r0
  474=>x"0EDB",	-- 0000111011011011  sbc	r3, r3, r3
  475=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  476=>x"08C9",	-- 0000100011001001  add	r1, r1, r3
  477=>x"0D00",	-- 0000110100000000  adc	r0, r0, r4
  478=>x"062D",	-- 0000011000101101  dec	r5, r5
  479=>x"BE6C",	-- 1011111001101100  brine	r5, mult_16_16.loop
  480=>x"E383",	-- 1110001110000011  ba	-, r6
  481=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  482=>x"C084",	-- 1100000010000100  li	r4, 16
  483=>x"0800",	-- 0000100000000000  add	r0, r0, r0
  484=>x"0C49",	-- 0000110001001001  adc	r1, r1, r1
  485=>x"0A8B",	-- 0000101010001011  sub	r3, r1, r2
  486=>x"80DD",	-- 1000000011011101  brilt	r3, div_16_16.skip
  487=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  488=>x"0400",	-- 0000010000000000  inc	r0, r0
  489=>x"0624",	-- 0000011000100100  dec	r4, r4
  490=>x"BE64",	-- 1011111001100100  brine	r4, div_16_16.loop
  491=>x"E383",	-- 1110001110000011  ba	-, r6
  492=>x"2400",	-- 0010010000000000  xor	r0, r0, r0
  493=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  494=>x"8250",	-- 1000001001010000  brieq	r2, fact_16.end
  495=>x"0409",	-- 0000010000001001  inc	r1, r1
  496=>x"1008",	-- 0001000000001000  mova	r0, r1
  497=>x"FAC6",	-- 1111101011000110  bail	-, r6, mult_16_16
  498=>x"01D5",	-- 0000000111010101  
  499=>x"8104",	-- 1000000100000100  brine	r0, fact_16.overflow
  500=>x"01D5",	-- 0000000111010101  
  501=>x"0612",	-- 0000011000010010  dec	r2, r2
  502=>x"BE94",	-- 1011111010010100  brine	r2, fact_16.loop
  503=>x"E383",	-- 1110001110000011  ba	-, r6
  504=>x"063F",	-- 0000011000111111  dec	r7, r7
  505=>x"D23E",	-- 1101001000111110  sw	r6, r7
  506=>x"D013",	-- 1101000000010011  lw	r3, r2
  507=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  508=>x"84D8",	-- 1000010011011000  brieq	r3, puts.end
  509=>x"063F",	-- 0000011000111111  dec	r7, r7
  510=>x"D23A",	-- 1101001000111010  sw	r2, r7
  511=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  512=>x"0212",	-- 0000001000010010  
  513=>x"D03A",	-- 1101000000111010  lw	r2, r7
  514=>x"043F",	-- 0000010000111111  inc	r7, r7
  515=>x"D013",	-- 1101000000010011  lw	r3, r2
  516=>x"4E1B",	-- 0100111000011011  shl	r3, r3, 7
  517=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  518=>x"8258",	-- 1000001001011000  brieq	r3, puts.end
  519=>x"063F",	-- 0000011000111111  dec	r7, r7
  520=>x"D23A",	-- 1101001000111010  sw	r2, r7
  521=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  522=>x"0212",	-- 0000001000010010  
  523=>x"D03A",	-- 1101000000111010  lw	r2, r7
  524=>x"043F",	-- 0000010000111111  inc	r7, r7
  525=>x"0412",	-- 0000010000010010  inc	r2, r2
  526=>x"BB03",	-- 1011101100000011  bri	-, puts.loop
  527=>x"D03E",	-- 1101000000111110  lw	r6, r7
  528=>x"043F",	-- 0000010000111111  inc	r7, r7
  529=>x"E383",	-- 1110001110000011  ba	-, r6
  530=>x"063F",	-- 0000011000111111  dec	r7, r7
  531=>x"D23E",	-- 1101001000111110  sw	r6, r7
  532=>x"063F",	-- 0000011000111111  dec	r7, r7
  533=>x"D238",	-- 1101001000111000  sw	r0, r7
  534=>x"063F",	-- 0000011000111111  dec	r7, r7
  535=>x"D239",	-- 1101001000111001  sw	r1, r7
  536=>x"FFF2",	-- 1111111111110010  liw	r2, font_map
  537=>x"12C0",	-- 0001001011000000  
  538=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  539=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  540=>x"C043",	-- 1100000001000011  li	r3, 8
  541=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  542=>x"025D",	-- 0000001001011101  
  543=>x"D039",	-- 1101000000111001  lw	r1, r7
  544=>x"043F",	-- 0000010000111111  inc	r7, r7
  545=>x"D038",	-- 1101000000111000  lw	r0, r7
  546=>x"043F",	-- 0000010000111111  inc	r7, r7
  547=>x"0400",	-- 0000010000000000  inc	r0, r0
  548=>x"D03E",	-- 1101000000111110  lw	r6, r7
  549=>x"043F",	-- 0000010000111111  inc	r7, r7
  550=>x"E383",	-- 1110001110000011  ba	-, r6
  551=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  552=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  553=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  554=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  555=>x"C0A0",	-- 1100000010100000  li	r0, 20
  556=>x"D011",	-- 1101000000010001  lw	r1, r2
  557=>x"D221",	-- 1101001000100001  sw	r1, r4
  558=>x"0412",	-- 0000010000010010  inc	r2, r2
  559=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  560=>x"061B",	-- 0000011000011011  dec	r3, r3
  561=>x"BEDC",	-- 1011111011011100  brine	r3, put_sprite_16_aligned.loop
  562=>x"E383",	-- 1110001110000011  ba	-, r6
  563=>x"C07D",	-- 1100000001111101  li	r5, 15
  564=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  565=>x"6600",	-- 0110011000000000  shr	r0, r0, 3
  566=>x"BC68",	-- 1011110001101000  brieq	r5, put_sprite_16_aligned
  567=>x"062D",	-- 0000011000101101  dec	r5, r5
  568=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  569=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  570=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  571=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  572=>x"063F",	-- 0000011000111111  dec	r7, r7
  573=>x"D23B",	-- 1101001000111011  sw	r3, r7
  574=>x"D011",	-- 1101000000010001  lw	r1, r2
  575=>x"CFF8",	-- 1100111111111000  li	r0, -1
  576=>x"3D40",	-- 0011110101000000  rsr	r0, r0, r5
  577=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  578=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  579=>x"D023",	-- 1101000000100011  lw	r3, r4
  580=>x"2600",	-- 0010011000000000  not	r0, r0
  581=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  582=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  583=>x"D221",	-- 1101001000100001  sw	r1, r4
  584=>x"0424",	-- 0000010000100100  inc	r4, r4
  585=>x"D011",	-- 1101000000010001  lw	r1, r2
  586=>x"262D",	-- 0010011000101101  not	r5, r5
  587=>x"CFF8",	-- 1100111111111000  li	r0, -1
  588=>x"3F40",	-- 0011111101000000  rsl	r0, r0, r5
  589=>x"3B49",	-- 0011101101001001  rrl	r1, r1, r5
  590=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  591=>x"262D",	-- 0010011000101101  not	r5, r5
  592=>x"D023",	-- 1101000000100011  lw	r3, r4
  593=>x"2600",	-- 0010011000000000  not	r0, r0
  594=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  595=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  596=>x"D221",	-- 1101001000100001  sw	r1, r4
  597=>x"0412",	-- 0000010000010010  inc	r2, r2
  598=>x"C098",	-- 1100000010011000  li	r0, 19
  599=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  600=>x"D03B",	-- 1101000000111011  lw	r3, r7
  601=>x"043F",	-- 0000010000111111  inc	r7, r7
  602=>x"061B",	-- 0000011000011011  dec	r3, r3
  603=>x"B85C",	-- 1011100001011100  brine	r3, put_sprite_16.loop
  604=>x"E383",	-- 1110001110000011  ba	-, r6
  605=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  606=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  607=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  608=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  609=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  610=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  611=>x"C0A5",	-- 1100000010100101  li	r5, 20
  612=>x"8404",	-- 1000010000000100  brine	r0, put_sprite_8_aligned.loop1
  613=>x"D010",	-- 1101000000010000  lw	r0, r2
  614=>x"D021",	-- 1101000000100001  lw	r1, r4
  615=>x"1A41",	-- 0001101001000001  mixhl	r1, r0, r1
  616=>x"D221",	-- 1101001000100001  sw	r1, r4
  617=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  618=>x"061B",	-- 0000011000011011  dec	r3, r3
  619=>x"E398",	-- 1110001110011000  baeq	r3, r6
  620=>x"D021",	-- 1101000000100001  lw	r1, r4
  621=>x"1E41",	-- 0001111001000001  mixll	r1, r0, r1
  622=>x"D221",	-- 1101001000100001  sw	r1, r4
  623=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  624=>x"0412",	-- 0000010000010010  inc	r2, r2
  625=>x"061B",	-- 0000011000011011  dec	r3, r3
  626=>x"E398",	-- 1110001110011000  baeq	r3, r6
  627=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop0
  628=>x"D010",	-- 1101000000010000  lw	r0, r2
  629=>x"D021",	-- 1101000000100001  lw	r1, r4
  630=>x"1809",	-- 0001100000001001  mixhh	r1, r1, r0
  631=>x"D221",	-- 1101001000100001  sw	r1, r4
  632=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  633=>x"061B",	-- 0000011000011011  dec	r3, r3
  634=>x"E398",	-- 1110001110011000  baeq	r3, r6
  635=>x"D021",	-- 1101000000100001  lw	r1, r4
  636=>x"1A09",	-- 0001101000001001  mixhl	r1, r1, r0
  637=>x"D221",	-- 1101001000100001  sw	r1, r4
  638=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  639=>x"0412",	-- 0000010000010010  inc	r2, r2
  640=>x"061B",	-- 0000011000011011  dec	r3, r3
  641=>x"E398",	-- 1110001110011000  baeq	r3, r6
  642=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop1
  643=>x"C03D",	-- 1100000000111101  li	r5, 7
  644=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  645=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  646=>x"B5E8",	-- 1011010111101000  brieq	r5, put_sprite_8_aligned
  647=>x"062D",	-- 0000011000101101  dec	r5, r5
  648=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  649=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  650=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  651=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  652=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  653=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  654=>x"8A04",	-- 1000101000000100  brine	r0, put_sprite_8.loop1
  655=>x"D010",	-- 1101000000010000  lw	r0, r2
  656=>x"063F",	-- 0000011000111111  dec	r7, r7
  657=>x"D23A",	-- 1101001000111010  sw	r2, r7
  658=>x"C802",	-- 1100100000000010  li	r2, 0x100
  659=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  660=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  661=>x"D021",	-- 1101000000100001  lw	r1, r4
  662=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  663=>x"2612",	-- 0010011000010010  not	r2, r2
  664=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  665=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  666=>x"D221",	-- 1101001000100001  sw	r1, r4
  667=>x"C0A1",	-- 1100000010100001  li	r1, 20
  668=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  669=>x"D03A",	-- 1101000000111010  lw	r2, r7
  670=>x"043F",	-- 0000010000111111  inc	r7, r7
  671=>x"061B",	-- 0000011000011011  dec	r3, r3
  672=>x"E398",	-- 1110001110011000  baeq	r3, r6
  673=>x"D010",	-- 1101000000010000  lw	r0, r2
  674=>x"063F",	-- 0000011000111111  dec	r7, r7
  675=>x"D23A",	-- 1101001000111010  sw	r2, r7
  676=>x"1E00",	-- 0001111000000000  mixll	r0, r0, r0
  677=>x"C802",	-- 1100100000000010  li	r2, 0x100
  678=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  679=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  680=>x"D021",	-- 1101000000100001  lw	r1, r4
  681=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  682=>x"2612",	-- 0010011000010010  not	r2, r2
  683=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  684=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  685=>x"D221",	-- 1101001000100001  sw	r1, r4
  686=>x"C0A1",	-- 1100000010100001  li	r1, 20
  687=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  688=>x"D03A",	-- 1101000000111010  lw	r2, r7
  689=>x"043F",	-- 0000010000111111  inc	r7, r7
  690=>x"0412",	-- 0000010000010010  inc	r2, r2
  691=>x"061B",	-- 0000011000011011  dec	r3, r3
  692=>x"E398",	-- 1110001110011000  baeq	r3, r6
  693=>x"B683",	-- 1011011010000011  bri	-, put_sprite_8.loop0
  694=>x"D010",	-- 1101000000010000  lw	r0, r2
  695=>x"063F",	-- 0000011000111111  dec	r7, r7
  696=>x"D23A",	-- 1101001000111010  sw	r2, r7
  697=>x"063F",	-- 0000011000111111  dec	r7, r7
  698=>x"D23B",	-- 1101001000111011  sw	r3, r7
  699=>x"C802",	-- 1100100000000010  li	r2, 0x100
  700=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  701=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  702=>x"2080",	-- 0010000010000000  and	r0, r0, r2
  703=>x"D021",	-- 1101000000100001  lw	r1, r4
  704=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
  705=>x"261B",	-- 0010011000011011  not	r3, r3
  706=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  707=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
  708=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  709=>x"D221",	-- 1101001000100001  sw	r1, r4
  710=>x"0424",	-- 0000010000100100  inc	r4, r4
  711=>x"D021",	-- 1101000000100001  lw	r1, r4
  712=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  713=>x"261B",	-- 0010011000011011  not	r3, r3
  714=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  715=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
  716=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  717=>x"D221",	-- 1101001000100001  sw	r1, r4
  718=>x"C099",	-- 1100000010011001  li	r1, 19
  719=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  720=>x"D03B",	-- 1101000000111011  lw	r3, r7
  721=>x"043F",	-- 0000010000111111  inc	r7, r7
  722=>x"D03A",	-- 1101000000111010  lw	r2, r7
  723=>x"043F",	-- 0000010000111111  inc	r7, r7
  724=>x"061B",	-- 0000011000011011  dec	r3, r3
  725=>x"E398",	-- 1110001110011000  baeq	r3, r6
  726=>x"D010",	-- 1101000000010000  lw	r0, r2
  727=>x"4E00",	-- 0100111000000000  shl	r0, r0, 7
  728=>x"063F",	-- 0000011000111111  dec	r7, r7
  729=>x"D23A",	-- 1101001000111010  sw	r2, r7
  730=>x"063F",	-- 0000011000111111  dec	r7, r7
  731=>x"D23B",	-- 1101001000111011  sw	r3, r7
  732=>x"C802",	-- 1100100000000010  li	r2, 0x100
  733=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  734=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  735=>x"2080",	-- 0010000010000000  and	r0, r0, r2
  736=>x"D021",	-- 1101000000100001  lw	r1, r4
  737=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
  738=>x"261B",	-- 0010011000011011  not	r3, r3
  739=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  740=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
  741=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  742=>x"D221",	-- 1101001000100001  sw	r1, r4
  743=>x"0424",	-- 0000010000100100  inc	r4, r4
  744=>x"D021",	-- 1101000000100001  lw	r1, r4
  745=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  746=>x"261B",	-- 0010011000011011  not	r3, r3
  747=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  748=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
  749=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  750=>x"D221",	-- 1101001000100001  sw	r1, r4
  751=>x"C099",	-- 1100000010011001  li	r1, 19
  752=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  753=>x"D03B",	-- 1101000000111011  lw	r3, r7
  754=>x"043F",	-- 0000010000111111  inc	r7, r7
  755=>x"D03A",	-- 1101000000111010  lw	r2, r7
  756=>x"043F",	-- 0000010000111111  inc	r7, r7
  757=>x"0412",	-- 0000010000010010  inc	r2, r2
  758=>x"061B",	-- 0000011000011011  dec	r3, r3
  759=>x"E398",	-- 1110001110011000  baeq	r3, r6
  760=>x"AF83",	-- 1010111110000011  bri	-, put_sprite_8.loop1
    others => x"0000"
    );
begin
  process(CLK)
  begin
    if (CLK'event AND CLK='1') then
      D <= m(to_integer(unsigned(AD)));
    end if;
  end process;
end Behavioral;
