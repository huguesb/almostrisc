library ieee;
use ieee.std_logic_1164.ALL;
use ieee.numeric_std.ALL;
library UNISIM;
use UNISIM.Vcomponents.ALL;
use work.dram_data_pkg.all;

entity RAMDoublePort is
   port ( AD1 : in  STD_LOGIC_VECTOR (12 downto 0);
          AD2 : in  STD_LOGIC_VECTOR (12 downto 0);
          DIN1 : in  STD_LOGIC_VECTOR (15 downto 0);
          DOUT1 : out  STD_LOGIC_VECTOR (15 downto 0);
          WE1 : in  STD_LOGIC;
          DOUT2 : out  STD_LOGIC_VECTOR (15 downto 0);
          OE1 : in  STD_LOGIC;
          CE1 : in  STD_LOGIC;
          CLK : in STD_LOGIC
    );
end RAMDoublePort;

architecture BEHAVIORAL of RAMDoublePort is
	component RAMB16_S9_S9
		generic
		(
			INIT_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_0A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_0B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_0C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_0D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_0E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_0F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INITP_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INITP_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INITP_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INITP_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INITP_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INITP_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INITP_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INITP_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_A : bit_vector := X"000";
			INIT_B : bit_vector := X"000";
			SIM_COLLISION_CHECK : string := "ALL";
			SRVAL_A : bit_vector := X"000";
			SRVAL_B : bit_vector := X"000";
			WRITE_MODE_A : string := "WRITE_FIRST";
			WRITE_MODE_B : string := "READ_FIRST"
		);
		port
		(
			DOA : out std_logic_vector(7 downto 0);
			DOB : out std_logic_vector(7 downto 0);
			DOPA : out std_logic_vector(0 downto 0);
			DOPB : out std_logic_vector(0 downto 0);
			ADDRA : in std_logic_vector(10 downto 0);
			ADDRB : in std_logic_vector(10 downto 0);
			CLKA : in std_ulogic;
			CLKB : in std_ulogic;
			DIA : in std_logic_vector(7 downto 0);
			DIB : in std_logic_vector(7 downto 0);
			DIPA : in std_logic_vector(0 downto 0);
			DIPB : in std_logic_vector(0 downto 0);
			ENA : in std_ulogic;
			ENB : in std_ulogic;
			SSRA : in std_ulogic;
			SSRB : in std_ulogic;
			WEA : in std_ulogic;
			WEB : in std_ulogic
		);
	end component;
	
	type vmb is array (3 downto 0) of std_logic_vector(15 downto 0);
	signal douta, doutb : vmb;
	signal phigh, plow : std_logic;
	signal pout : std_logic_vector(15 downto 0);
begin
	plow <= ((DIN1(7) xor DIN1(6)) xor (DIN1(5) xor DIN1(4))) xor ((DIN1(3) xor DIN1(2)) xor (DIN1(1) xor DIN1(0)));
	phigh <= ((DIN1(15) xor DIN1(14)) xor (DIN1(13) xor DIN1(12))) xor ((DIN1(11) xor DIN1(10)) xor (DIN1(9) xor DIN1(8)));
	
	XLXI_0 : RAMB16_S9_S9
	generic map (
		INIT_00=>cRAMDoublePort_XLXI_0_INIT_00,
		INIT_01=>cRAMDoublePort_XLXI_0_INIT_01,
		INIT_02=>cRAMDoublePort_XLXI_0_INIT_02,
		INIT_03=>cRAMDoublePort_XLXI_0_INIT_03,
		INIT_04=>cRAMDoublePort_XLXI_0_INIT_04,
		INIT_05=>cRAMDoublePort_XLXI_0_INIT_05,
		INIT_06=>cRAMDoublePort_XLXI_0_INIT_06,
		INIT_07=>cRAMDoublePort_XLXI_0_INIT_07,
		INIT_08=>cRAMDoublePort_XLXI_0_INIT_08,
		INIT_09=>cRAMDoublePort_XLXI_0_INIT_09,
		INIT_0a=>cRAMDoublePort_XLXI_0_INIT_0A,
		INIT_0b=>cRAMDoublePort_XLXI_0_INIT_0B,
		INIT_0c=>cRAMDoublePort_XLXI_0_INIT_0C,
		INIT_0d=>cRAMDoublePort_XLXI_0_INIT_0D,
		INIT_0e=>cRAMDoublePort_XLXI_0_INIT_0E,
		INIT_0f=>cRAMDoublePort_XLXI_0_INIT_0F,
		INIT_10=>cRAMDoublePort_XLXI_0_INIT_10,
		INIT_11=>cRAMDoublePort_XLXI_0_INIT_11,
		INIT_12=>cRAMDoublePort_XLXI_0_INIT_12,
		INIT_13=>cRAMDoublePort_XLXI_0_INIT_13,
		INIT_14=>cRAMDoublePort_XLXI_0_INIT_14,
		INIT_15=>cRAMDoublePort_XLXI_0_INIT_15,
		INIT_16=>cRAMDoublePort_XLXI_0_INIT_16,
		INIT_17=>cRAMDoublePort_XLXI_0_INIT_17,
		INIT_18=>cRAMDoublePort_XLXI_0_INIT_18,
		INIT_19=>cRAMDoublePort_XLXI_0_INIT_19,
		INIT_1a=>cRAMDoublePort_XLXI_0_INIT_1A,
		INIT_1b=>cRAMDoublePort_XLXI_0_INIT_1B,
		INIT_1c=>cRAMDoublePort_XLXI_0_INIT_1C,
		INIT_1d=>cRAMDoublePort_XLXI_0_INIT_1D,
		INIT_1e=>cRAMDoublePort_XLXI_0_INIT_1E,
		INIT_1f=>cRAMDoublePort_XLXI_0_INIT_1F,
		INIT_20=>cRAMDoublePort_XLXI_0_INIT_20,
		INIT_21=>cRAMDoublePort_XLXI_0_INIT_21,
		INIT_22=>cRAMDoublePort_XLXI_0_INIT_22,
		INIT_23=>cRAMDoublePort_XLXI_0_INIT_23,
		INIT_24=>cRAMDoublePort_XLXI_0_INIT_24,
		INIT_25=>cRAMDoublePort_XLXI_0_INIT_25,
		INIT_26=>cRAMDoublePort_XLXI_0_INIT_26,
		INIT_27=>cRAMDoublePort_XLXI_0_INIT_27,
		INIT_28=>cRAMDoublePort_XLXI_0_INIT_28,
		INIT_29=>cRAMDoublePort_XLXI_0_INIT_29,
		INIT_2a=>cRAMDoublePort_XLXI_0_INIT_2A,
		INIT_2b=>cRAMDoublePort_XLXI_0_INIT_2B,
		INIT_2c=>cRAMDoublePort_XLXI_0_INIT_2C,
		INIT_2d=>cRAMDoublePort_XLXI_0_INIT_2D,
		INIT_2e=>cRAMDoublePort_XLXI_0_INIT_2E,
		INIT_2f=>cRAMDoublePort_XLXI_0_INIT_2F,
		INIT_30=>cRAMDoublePort_XLXI_0_INIT_30,
		INIT_31=>cRAMDoublePort_XLXI_0_INIT_31,
		INIT_32=>cRAMDoublePort_XLXI_0_INIT_32,
		INIT_33=>cRAMDoublePort_XLXI_0_INIT_33,
		INIT_34=>cRAMDoublePort_XLXI_0_INIT_34,
		INIT_35=>cRAMDoublePort_XLXI_0_INIT_35,
		INIT_36=>cRAMDoublePort_XLXI_0_INIT_36,
		INIT_37=>cRAMDoublePort_XLXI_0_INIT_37,
		INIT_38=>cRAMDoublePort_XLXI_0_INIT_38,
		INIT_39=>cRAMDoublePort_XLXI_0_INIT_39,
		INIT_3a=>cRAMDoublePort_XLXI_0_INIT_3A,
		INIT_3b=>cRAMDoublePort_XLXI_0_INIT_3B,
		INIT_3c=>cRAMDoublePort_XLXI_0_INIT_3C,
		INIT_3d=>cRAMDoublePort_XLXI_0_INIT_3D,
		INIT_3e=>cRAMDoublePort_XLXI_0_INIT_3E,
		INIT_3f=>cRAMDoublePort_XLXI_0_INIT_3F
	)
	port map (
		CLKA=>CLK,
		ENA=>CE1,
		WEA=>WE1,
		SSRA=>'0',
		ADDRA=>AD1(10 downto 0),
		DIA=>DIN1(7 downto 0),
		DIPA(0)=>plow,
		DOA=>douta(0)(7 downto 0),
		DOPA(0)=>pout(0),
		
		CLKB=>CLK,
		ENB=>'1',
		WEB=>'0',
		SSRB=>'0',
		ADDRB=>AD2(10 downto 0),
		DIB=>(others=>'0'),
		DIPB(0)=>'0',
		DOB=>doutb(0)(7 downto 0),
		DOPB(0)=>pout(1)
	);
	
	XLXI_1 : RAMB16_S9_S9
	generic map (
		INIT_00=>cRAMDoublePort_XLXI_1_INIT_00,
		INIT_01=>cRAMDoublePort_XLXI_1_INIT_01,
		INIT_02=>cRAMDoublePort_XLXI_1_INIT_02,
		INIT_03=>cRAMDoublePort_XLXI_1_INIT_03,
		INIT_04=>cRAMDoublePort_XLXI_1_INIT_04,
		INIT_05=>cRAMDoublePort_XLXI_1_INIT_05,
		INIT_06=>cRAMDoublePort_XLXI_1_INIT_06,
		INIT_07=>cRAMDoublePort_XLXI_1_INIT_07,
		INIT_08=>cRAMDoublePort_XLXI_1_INIT_08,
		INIT_09=>cRAMDoublePort_XLXI_1_INIT_09,
		INIT_0a=>cRAMDoublePort_XLXI_1_INIT_0A,
		INIT_0b=>cRAMDoublePort_XLXI_1_INIT_0B,
		INIT_0c=>cRAMDoublePort_XLXI_1_INIT_0C,
		INIT_0d=>cRAMDoublePort_XLXI_1_INIT_0D,
		INIT_0e=>cRAMDoublePort_XLXI_1_INIT_0E,
		INIT_0f=>cRAMDoublePort_XLXI_1_INIT_0F,
		INIT_10=>cRAMDoublePort_XLXI_1_INIT_10,
		INIT_11=>cRAMDoublePort_XLXI_1_INIT_11,
		INIT_12=>cRAMDoublePort_XLXI_1_INIT_12,
		INIT_13=>cRAMDoublePort_XLXI_1_INIT_13,
		INIT_14=>cRAMDoublePort_XLXI_1_INIT_14,
		INIT_15=>cRAMDoublePort_XLXI_1_INIT_15,
		INIT_16=>cRAMDoublePort_XLXI_1_INIT_16,
		INIT_17=>cRAMDoublePort_XLXI_1_INIT_17,
		INIT_18=>cRAMDoublePort_XLXI_1_INIT_18,
		INIT_19=>cRAMDoublePort_XLXI_1_INIT_19,
		INIT_1a=>cRAMDoublePort_XLXI_1_INIT_1A,
		INIT_1b=>cRAMDoublePort_XLXI_1_INIT_1B,
		INIT_1c=>cRAMDoublePort_XLXI_1_INIT_1C,
		INIT_1d=>cRAMDoublePort_XLXI_1_INIT_1D,
		INIT_1e=>cRAMDoublePort_XLXI_1_INIT_1E,
		INIT_1f=>cRAMDoublePort_XLXI_1_INIT_1F,
		INIT_20=>cRAMDoublePort_XLXI_1_INIT_20,
		INIT_21=>cRAMDoublePort_XLXI_1_INIT_21,
		INIT_22=>cRAMDoublePort_XLXI_1_INIT_22,
		INIT_23=>cRAMDoublePort_XLXI_1_INIT_23,
		INIT_24=>cRAMDoublePort_XLXI_1_INIT_24,
		INIT_25=>cRAMDoublePort_XLXI_1_INIT_25,
		INIT_26=>cRAMDoublePort_XLXI_1_INIT_26,
		INIT_27=>cRAMDoublePort_XLXI_1_INIT_27,
		INIT_28=>cRAMDoublePort_XLXI_1_INIT_28,
		INIT_29=>cRAMDoublePort_XLXI_1_INIT_29,
		INIT_2a=>cRAMDoublePort_XLXI_1_INIT_2A,
		INIT_2b=>cRAMDoublePort_XLXI_1_INIT_2B,
		INIT_2c=>cRAMDoublePort_XLXI_1_INIT_2C,
		INIT_2d=>cRAMDoublePort_XLXI_1_INIT_2D,
		INIT_2e=>cRAMDoublePort_XLXI_1_INIT_2E,
		INIT_2f=>cRAMDoublePort_XLXI_1_INIT_2F,
		INIT_30=>cRAMDoublePort_XLXI_1_INIT_30,
		INIT_31=>cRAMDoublePort_XLXI_1_INIT_31,
		INIT_32=>cRAMDoublePort_XLXI_1_INIT_32,
		INIT_33=>cRAMDoublePort_XLXI_1_INIT_33,
		INIT_34=>cRAMDoublePort_XLXI_1_INIT_34,
		INIT_35=>cRAMDoublePort_XLXI_1_INIT_35,
		INIT_36=>cRAMDoublePort_XLXI_1_INIT_36,
		INIT_37=>cRAMDoublePort_XLXI_1_INIT_37,
		INIT_38=>cRAMDoublePort_XLXI_1_INIT_38,
		INIT_39=>cRAMDoublePort_XLXI_1_INIT_39,
		INIT_3a=>cRAMDoublePort_XLXI_1_INIT_3A,
		INIT_3b=>cRAMDoublePort_XLXI_1_INIT_3B,
		INIT_3c=>cRAMDoublePort_XLXI_1_INIT_3C,
		INIT_3d=>cRAMDoublePort_XLXI_1_INIT_3D,
		INIT_3e=>cRAMDoublePort_XLXI_1_INIT_3E,
		INIT_3f=>cRAMDoublePort_XLXI_1_INIT_3F
	)
	port map (
		CLKA=>CLK,
		ENA=>CE1,
		WEA=>WE1,
		SSRA=>'0',
		ADDRA=>AD1(10 downto 0),
		DIA=>DIN1(7 downto 0),
		DIPA(0)=>phigh,
		DOA=>douta(0)(15 downto 8),
		DOPA(0)=>pout(2),
		
		CLKB=>CLK,
		ENB=>'1',
		WEB=>'0',
		SSRB=>'0',
		ADDRB=>AD2(10 downto 0),
		DIB=>(others=>'0'),
		DIPB(0)=>'0',
		DOB=>doutb(0)(15 downto 8),
		DOPB(0)=>pout(3)
	);
	
	XLXI_2 : RAMB16_S9_S9
	generic map (
		INIT_00=>cRAMDoublePort_XLXI_2_INIT_00,
		INIT_01=>cRAMDoublePort_XLXI_2_INIT_01,
		INIT_02=>cRAMDoublePort_XLXI_2_INIT_02,
		INIT_03=>cRAMDoublePort_XLXI_2_INIT_03,
		INIT_04=>cRAMDoublePort_XLXI_2_INIT_04,
		INIT_05=>cRAMDoublePort_XLXI_2_INIT_05,
		INIT_06=>cRAMDoublePort_XLXI_2_INIT_06,
		INIT_07=>cRAMDoublePort_XLXI_2_INIT_07,
		INIT_08=>cRAMDoublePort_XLXI_2_INIT_08,
		INIT_09=>cRAMDoublePort_XLXI_2_INIT_09,
		INIT_0a=>cRAMDoublePort_XLXI_2_INIT_0A,
		INIT_0b=>cRAMDoublePort_XLXI_2_INIT_0B,
		INIT_0c=>cRAMDoublePort_XLXI_2_INIT_0C,
		INIT_0d=>cRAMDoublePort_XLXI_2_INIT_0D,
		INIT_0e=>cRAMDoublePort_XLXI_2_INIT_0E,
		INIT_0f=>cRAMDoublePort_XLXI_2_INIT_0F,
		INIT_10=>cRAMDoublePort_XLXI_2_INIT_10,
		INIT_11=>cRAMDoublePort_XLXI_2_INIT_11,
		INIT_12=>cRAMDoublePort_XLXI_2_INIT_12,
		INIT_13=>cRAMDoublePort_XLXI_2_INIT_13,
		INIT_14=>cRAMDoublePort_XLXI_2_INIT_14,
		INIT_15=>cRAMDoublePort_XLXI_2_INIT_15,
		INIT_16=>cRAMDoublePort_XLXI_2_INIT_16,
		INIT_17=>cRAMDoublePort_XLXI_2_INIT_17,
		INIT_18=>cRAMDoublePort_XLXI_2_INIT_18,
		INIT_19=>cRAMDoublePort_XLXI_2_INIT_19,
		INIT_1a=>cRAMDoublePort_XLXI_2_INIT_1A,
		INIT_1b=>cRAMDoublePort_XLXI_2_INIT_1B,
		INIT_1c=>cRAMDoublePort_XLXI_2_INIT_1C,
		INIT_1d=>cRAMDoublePort_XLXI_2_INIT_1D,
		INIT_1e=>cRAMDoublePort_XLXI_2_INIT_1E,
		INIT_1f=>cRAMDoublePort_XLXI_2_INIT_1F,
		INIT_20=>cRAMDoublePort_XLXI_2_INIT_20,
		INIT_21=>cRAMDoublePort_XLXI_2_INIT_21,
		INIT_22=>cRAMDoublePort_XLXI_2_INIT_22,
		INIT_23=>cRAMDoublePort_XLXI_2_INIT_23,
		INIT_24=>cRAMDoublePort_XLXI_2_INIT_24,
		INIT_25=>cRAMDoublePort_XLXI_2_INIT_25,
		INIT_26=>cRAMDoublePort_XLXI_2_INIT_26,
		INIT_27=>cRAMDoublePort_XLXI_2_INIT_27,
		INIT_28=>cRAMDoublePort_XLXI_2_INIT_28,
		INIT_29=>cRAMDoublePort_XLXI_2_INIT_29,
		INIT_2a=>cRAMDoublePort_XLXI_2_INIT_2A,
		INIT_2b=>cRAMDoublePort_XLXI_2_INIT_2B,
		INIT_2c=>cRAMDoublePort_XLXI_2_INIT_2C,
		INIT_2d=>cRAMDoublePort_XLXI_2_INIT_2D,
		INIT_2e=>cRAMDoublePort_XLXI_2_INIT_2E,
		INIT_2f=>cRAMDoublePort_XLXI_2_INIT_2F,
		INIT_30=>cRAMDoublePort_XLXI_2_INIT_30,
		INIT_31=>cRAMDoublePort_XLXI_2_INIT_31,
		INIT_32=>cRAMDoublePort_XLXI_2_INIT_32,
		INIT_33=>cRAMDoublePort_XLXI_2_INIT_33,
		INIT_34=>cRAMDoublePort_XLXI_2_INIT_34,
		INIT_35=>cRAMDoublePort_XLXI_2_INIT_35,
		INIT_36=>cRAMDoublePort_XLXI_2_INIT_36,
		INIT_37=>cRAMDoublePort_XLXI_2_INIT_37,
		INIT_38=>cRAMDoublePort_XLXI_2_INIT_38,
		INIT_39=>cRAMDoublePort_XLXI_2_INIT_39,
		INIT_3a=>cRAMDoublePort_XLXI_2_INIT_3A,
		INIT_3b=>cRAMDoublePort_XLXI_2_INIT_3B,
		INIT_3c=>cRAMDoublePort_XLXI_2_INIT_3C,
		INIT_3d=>cRAMDoublePort_XLXI_2_INIT_3D,
		INIT_3e=>cRAMDoublePort_XLXI_2_INIT_3E,
		INIT_3f=>cRAMDoublePort_XLXI_2_INIT_3F
	)
	port map (
		CLKA=>CLK,
		ENA=>CE1,
		WEA=>WE1,
		SSRA=>'0',
		ADDRA=>AD1(10 downto 0),
		DIA=>DIN1(7 downto 0),
		DIPA(0)=>plow,
		DOA=>douta(1)(7 downto 0),
		DOPA(0)=>pout(4),
		
		CLKB=>CLK,
		ENB=>'1',
		WEB=>'0',
		SSRB=>'0',
		ADDRB=>AD2(10 downto 0),
		DIB=>(others=>'0'),
		DIPB(0)=>'0',
		DOB=>doutb(1)(7 downto 0),
		DOPB(0)=>pout(5)
	);
	
	XLXI_3 : RAMB16_S9_S9
	generic map (
		INIT_00=>cRAMDoublePort_XLXI_3_INIT_00,
		INIT_01=>cRAMDoublePort_XLXI_3_INIT_01,
		INIT_02=>cRAMDoublePort_XLXI_3_INIT_02,
		INIT_03=>cRAMDoublePort_XLXI_3_INIT_03,
		INIT_04=>cRAMDoublePort_XLXI_3_INIT_04,
		INIT_05=>cRAMDoublePort_XLXI_3_INIT_05,
		INIT_06=>cRAMDoublePort_XLXI_3_INIT_06,
		INIT_07=>cRAMDoublePort_XLXI_3_INIT_07,
		INIT_08=>cRAMDoublePort_XLXI_3_INIT_08,
		INIT_09=>cRAMDoublePort_XLXI_3_INIT_09,
		INIT_0a=>cRAMDoublePort_XLXI_3_INIT_0A,
		INIT_0b=>cRAMDoublePort_XLXI_3_INIT_0B,
		INIT_0c=>cRAMDoublePort_XLXI_3_INIT_0C,
		INIT_0d=>cRAMDoublePort_XLXI_3_INIT_0D,
		INIT_0e=>cRAMDoublePort_XLXI_3_INIT_0E,
		INIT_0f=>cRAMDoublePort_XLXI_3_INIT_0F,
		INIT_10=>cRAMDoublePort_XLXI_3_INIT_10,
		INIT_11=>cRAMDoublePort_XLXI_3_INIT_11,
		INIT_12=>cRAMDoublePort_XLXI_3_INIT_12,
		INIT_13=>cRAMDoublePort_XLXI_3_INIT_13,
		INIT_14=>cRAMDoublePort_XLXI_3_INIT_14,
		INIT_15=>cRAMDoublePort_XLXI_3_INIT_15,
		INIT_16=>cRAMDoublePort_XLXI_3_INIT_16,
		INIT_17=>cRAMDoublePort_XLXI_3_INIT_17,
		INIT_18=>cRAMDoublePort_XLXI_3_INIT_18,
		INIT_19=>cRAMDoublePort_XLXI_3_INIT_19,
		INIT_1a=>cRAMDoublePort_XLXI_3_INIT_1A,
		INIT_1b=>cRAMDoublePort_XLXI_3_INIT_1B,
		INIT_1c=>cRAMDoublePort_XLXI_3_INIT_1C,
		INIT_1d=>cRAMDoublePort_XLXI_3_INIT_1D,
		INIT_1e=>cRAMDoublePort_XLXI_3_INIT_1E,
		INIT_1f=>cRAMDoublePort_XLXI_3_INIT_1F,
		INIT_20=>cRAMDoublePort_XLXI_3_INIT_20,
		INIT_21=>cRAMDoublePort_XLXI_3_INIT_21,
		INIT_22=>cRAMDoublePort_XLXI_3_INIT_22,
		INIT_23=>cRAMDoublePort_XLXI_3_INIT_23,
		INIT_24=>cRAMDoublePort_XLXI_3_INIT_24,
		INIT_25=>cRAMDoublePort_XLXI_3_INIT_25,
		INIT_26=>cRAMDoublePort_XLXI_3_INIT_26,
		INIT_27=>cRAMDoublePort_XLXI_3_INIT_27,
		INIT_28=>cRAMDoublePort_XLXI_3_INIT_28,
		INIT_29=>cRAMDoublePort_XLXI_3_INIT_29,
		INIT_2a=>cRAMDoublePort_XLXI_3_INIT_2A,
		INIT_2b=>cRAMDoublePort_XLXI_3_INIT_2B,
		INIT_2c=>cRAMDoublePort_XLXI_3_INIT_2C,
		INIT_2d=>cRAMDoublePort_XLXI_3_INIT_2D,
		INIT_2e=>cRAMDoublePort_XLXI_3_INIT_2E,
		INIT_2f=>cRAMDoublePort_XLXI_3_INIT_2F,
		INIT_30=>cRAMDoublePort_XLXI_3_INIT_30,
		INIT_31=>cRAMDoublePort_XLXI_3_INIT_31,
		INIT_32=>cRAMDoublePort_XLXI_3_INIT_32,
		INIT_33=>cRAMDoublePort_XLXI_3_INIT_33,
		INIT_34=>cRAMDoublePort_XLXI_3_INIT_34,
		INIT_35=>cRAMDoublePort_XLXI_3_INIT_35,
		INIT_36=>cRAMDoublePort_XLXI_3_INIT_36,
		INIT_37=>cRAMDoublePort_XLXI_3_INIT_37,
		INIT_38=>cRAMDoublePort_XLXI_3_INIT_38,
		INIT_39=>cRAMDoublePort_XLXI_3_INIT_39,
		INIT_3a=>cRAMDoublePort_XLXI_3_INIT_3A,
		INIT_3b=>cRAMDoublePort_XLXI_3_INIT_3B,
		INIT_3c=>cRAMDoublePort_XLXI_3_INIT_3C,
		INIT_3d=>cRAMDoublePort_XLXI_3_INIT_3D,
		INIT_3e=>cRAMDoublePort_XLXI_3_INIT_3E,
		INIT_3f=>cRAMDoublePort_XLXI_3_INIT_3F
	)
	port map (
		CLKA=>CLK,
		ENA=>CE1,
		WEA=>WE1,
		SSRA=>'0',
		ADDRA=>AD1(10 downto 0),
		DIA=>DIN1(15 downto 8),
		DIPA(0)=>phigh,
		DOA=>douta(1)(15 downto 8),
		DOPA(0)=>pout(6),
		
		CLKB=>CLK,
		ENB=>'1',
		WEB=>'0',
		SSRB=>'0',
		ADDRB=>AD2(10 downto 0),
		DIB=>(others=>'0'),
		DIPB(0)=>'0',
		DOB=>doutb(1)(15 downto 8),
		DOPB(0)=>pout(7)
	);
	
	XLXI_4 : RAMB16_S9_S9
	generic map (
		INIT_00=>cRAMDoublePort_XLXI_4_INIT_00,
		INIT_01=>cRAMDoublePort_XLXI_4_INIT_01,
		INIT_02=>cRAMDoublePort_XLXI_4_INIT_02,
		INIT_03=>cRAMDoublePort_XLXI_4_INIT_03,
		INIT_04=>cRAMDoublePort_XLXI_4_INIT_04,
		INIT_05=>cRAMDoublePort_XLXI_4_INIT_05,
		INIT_06=>cRAMDoublePort_XLXI_4_INIT_06,
		INIT_07=>cRAMDoublePort_XLXI_4_INIT_07,
		INIT_08=>cRAMDoublePort_XLXI_4_INIT_08,
		INIT_09=>cRAMDoublePort_XLXI_4_INIT_09,
		INIT_0a=>cRAMDoublePort_XLXI_4_INIT_0A,
		INIT_0b=>cRAMDoublePort_XLXI_4_INIT_0B,
		INIT_0c=>cRAMDoublePort_XLXI_4_INIT_0C,
		INIT_0d=>cRAMDoublePort_XLXI_4_INIT_0D,
		INIT_0e=>cRAMDoublePort_XLXI_4_INIT_0E,
		INIT_0f=>cRAMDoublePort_XLXI_4_INIT_0F,
		INIT_10=>cRAMDoublePort_XLXI_4_INIT_10,
		INIT_11=>cRAMDoublePort_XLXI_4_INIT_11,
		INIT_12=>cRAMDoublePort_XLXI_4_INIT_12,
		INIT_13=>cRAMDoublePort_XLXI_4_INIT_13,
		INIT_14=>cRAMDoublePort_XLXI_4_INIT_14,
		INIT_15=>cRAMDoublePort_XLXI_4_INIT_15,
		INIT_16=>cRAMDoublePort_XLXI_4_INIT_16,
		INIT_17=>cRAMDoublePort_XLXI_4_INIT_17,
		INIT_18=>cRAMDoublePort_XLXI_4_INIT_18,
		INIT_19=>cRAMDoublePort_XLXI_4_INIT_19,
		INIT_1a=>cRAMDoublePort_XLXI_4_INIT_1A,
		INIT_1b=>cRAMDoublePort_XLXI_4_INIT_1B,
		INIT_1c=>cRAMDoublePort_XLXI_4_INIT_1C,
		INIT_1d=>cRAMDoublePort_XLXI_4_INIT_1D,
		INIT_1e=>cRAMDoublePort_XLXI_4_INIT_1E,
		INIT_1f=>cRAMDoublePort_XLXI_4_INIT_1F,
		INIT_20=>cRAMDoublePort_XLXI_4_INIT_20,
		INIT_21=>cRAMDoublePort_XLXI_4_INIT_21,
		INIT_22=>cRAMDoublePort_XLXI_4_INIT_22,
		INIT_23=>cRAMDoublePort_XLXI_4_INIT_23,
		INIT_24=>cRAMDoublePort_XLXI_4_INIT_24,
		INIT_25=>cRAMDoublePort_XLXI_4_INIT_25,
		INIT_26=>cRAMDoublePort_XLXI_4_INIT_26,
		INIT_27=>cRAMDoublePort_XLXI_4_INIT_27,
		INIT_28=>cRAMDoublePort_XLXI_4_INIT_28,
		INIT_29=>cRAMDoublePort_XLXI_4_INIT_29,
		INIT_2a=>cRAMDoublePort_XLXI_4_INIT_2A,
		INIT_2b=>cRAMDoublePort_XLXI_4_INIT_2B,
		INIT_2c=>cRAMDoublePort_XLXI_4_INIT_2C,
		INIT_2d=>cRAMDoublePort_XLXI_4_INIT_2D,
		INIT_2e=>cRAMDoublePort_XLXI_4_INIT_2E,
		INIT_2f=>cRAMDoublePort_XLXI_4_INIT_2F,
		INIT_30=>cRAMDoublePort_XLXI_4_INIT_30,
		INIT_31=>cRAMDoublePort_XLXI_4_INIT_31,
		INIT_32=>cRAMDoublePort_XLXI_4_INIT_32,
		INIT_33=>cRAMDoublePort_XLXI_4_INIT_33,
		INIT_34=>cRAMDoublePort_XLXI_4_INIT_34,
		INIT_35=>cRAMDoublePort_XLXI_4_INIT_35,
		INIT_36=>cRAMDoublePort_XLXI_4_INIT_36,
		INIT_37=>cRAMDoublePort_XLXI_4_INIT_37,
		INIT_38=>cRAMDoublePort_XLXI_4_INIT_38,
		INIT_39=>cRAMDoublePort_XLXI_4_INIT_39,
		INIT_3a=>cRAMDoublePort_XLXI_4_INIT_3A,
		INIT_3b=>cRAMDoublePort_XLXI_4_INIT_3B,
		INIT_3c=>cRAMDoublePort_XLXI_4_INIT_3C,
		INIT_3d=>cRAMDoublePort_XLXI_4_INIT_3D,
		INIT_3e=>cRAMDoublePort_XLXI_4_INIT_3E,
		INIT_3f=>cRAMDoublePort_XLXI_4_INIT_3F
	)
	port map (
		CLKA=>CLK,
		ENA=>CE1,
		WEA=>WE1,
		SSRA=>'0',
		ADDRA=>AD1(10 downto 0),
		DIA=>DIN1(7 downto 0),
		DIPA(0)=>plow,
		DOA=>douta(2)(7 downto 0),
		DOPA(0)=>pout(8),
		
		CLKB=>CLK,
		ENB=>'1',
		WEB=>'0',
		SSRB=>'0',
		ADDRB=>AD2(10 downto 0),
		DIB=>(others=>'0'),
		DIPB(0)=>'0',
		DOB=>doutb(2)(7 downto 0),
		DOPB(0)=>pout(9)
	);
	
	XLXI_5 : RAMB16_S9_S9
	generic map (
		INIT_00=>cRAMDoublePort_XLXI_5_INIT_00,
		INIT_01=>cRAMDoublePort_XLXI_5_INIT_01,
		INIT_02=>cRAMDoublePort_XLXI_5_INIT_02,
		INIT_03=>cRAMDoublePort_XLXI_5_INIT_03,
		INIT_04=>cRAMDoublePort_XLXI_5_INIT_04,
		INIT_05=>cRAMDoublePort_XLXI_5_INIT_05,
		INIT_06=>cRAMDoublePort_XLXI_5_INIT_06,
		INIT_07=>cRAMDoublePort_XLXI_5_INIT_07,
		INIT_08=>cRAMDoublePort_XLXI_5_INIT_08,
		INIT_09=>cRAMDoublePort_XLXI_5_INIT_09,
		INIT_0a=>cRAMDoublePort_XLXI_5_INIT_0A,
		INIT_0b=>cRAMDoublePort_XLXI_5_INIT_0B,
		INIT_0c=>cRAMDoublePort_XLXI_5_INIT_0C,
		INIT_0d=>cRAMDoublePort_XLXI_5_INIT_0D,
		INIT_0e=>cRAMDoublePort_XLXI_5_INIT_0E,
		INIT_0f=>cRAMDoublePort_XLXI_5_INIT_0F,
		INIT_10=>cRAMDoublePort_XLXI_5_INIT_10,
		INIT_11=>cRAMDoublePort_XLXI_5_INIT_11,
		INIT_12=>cRAMDoublePort_XLXI_5_INIT_12,
		INIT_13=>cRAMDoublePort_XLXI_5_INIT_13,
		INIT_14=>cRAMDoublePort_XLXI_5_INIT_14,
		INIT_15=>cRAMDoublePort_XLXI_5_INIT_15,
		INIT_16=>cRAMDoublePort_XLXI_5_INIT_16,
		INIT_17=>cRAMDoublePort_XLXI_5_INIT_17,
		INIT_18=>cRAMDoublePort_XLXI_5_INIT_18,
		INIT_19=>cRAMDoublePort_XLXI_5_INIT_19,
		INIT_1a=>cRAMDoublePort_XLXI_5_INIT_1A,
		INIT_1b=>cRAMDoublePort_XLXI_5_INIT_1B,
		INIT_1c=>cRAMDoublePort_XLXI_5_INIT_1C,
		INIT_1d=>cRAMDoublePort_XLXI_5_INIT_1D,
		INIT_1e=>cRAMDoublePort_XLXI_5_INIT_1E,
		INIT_1f=>cRAMDoublePort_XLXI_5_INIT_1F,
		INIT_20=>cRAMDoublePort_XLXI_5_INIT_20,
		INIT_21=>cRAMDoublePort_XLXI_5_INIT_21,
		INIT_22=>cRAMDoublePort_XLXI_5_INIT_22,
		INIT_23=>cRAMDoublePort_XLXI_5_INIT_23,
		INIT_24=>cRAMDoublePort_XLXI_5_INIT_24,
		INIT_25=>cRAMDoublePort_XLXI_5_INIT_25,
		INIT_26=>cRAMDoublePort_XLXI_5_INIT_26,
		INIT_27=>cRAMDoublePort_XLXI_5_INIT_27,
		INIT_28=>cRAMDoublePort_XLXI_5_INIT_28,
		INIT_29=>cRAMDoublePort_XLXI_5_INIT_29,
		INIT_2a=>cRAMDoublePort_XLXI_5_INIT_2A,
		INIT_2b=>cRAMDoublePort_XLXI_5_INIT_2B,
		INIT_2c=>cRAMDoublePort_XLXI_5_INIT_2C,
		INIT_2d=>cRAMDoublePort_XLXI_5_INIT_2D,
		INIT_2e=>cRAMDoublePort_XLXI_5_INIT_2E,
		INIT_2f=>cRAMDoublePort_XLXI_5_INIT_2F,
		INIT_30=>cRAMDoublePort_XLXI_5_INIT_30,
		INIT_31=>cRAMDoublePort_XLXI_5_INIT_31,
		INIT_32=>cRAMDoublePort_XLXI_5_INIT_32,
		INIT_33=>cRAMDoublePort_XLXI_5_INIT_33,
		INIT_34=>cRAMDoublePort_XLXI_5_INIT_34,
		INIT_35=>cRAMDoublePort_XLXI_5_INIT_35,
		INIT_36=>cRAMDoublePort_XLXI_5_INIT_36,
		INIT_37=>cRAMDoublePort_XLXI_5_INIT_37,
		INIT_38=>cRAMDoublePort_XLXI_5_INIT_38,
		INIT_39=>cRAMDoublePort_XLXI_5_INIT_39,
		INIT_3a=>cRAMDoublePort_XLXI_5_INIT_3A,
		INIT_3b=>cRAMDoublePort_XLXI_5_INIT_3B,
		INIT_3c=>cRAMDoublePort_XLXI_5_INIT_3C,
		INIT_3d=>cRAMDoublePort_XLXI_5_INIT_3D,
		INIT_3e=>cRAMDoublePort_XLXI_5_INIT_3E,
		INIT_3f=>cRAMDoublePort_XLXI_5_INIT_3F
	)
	port map (
		CLKA=>CLK,
		ENA=>CE1,
		WEA=>WE1,
		SSRA=>'0',
		ADDRA=>AD1(10 downto 0),
		DIA=>DIN1(15 downto 8),
		DIPA(0)=>phigh,
		DOA=>douta(2)(15 downto 8),
		DOPA(0)=>pout(10),
		
		CLKB=>CLK,
		ENB=>'1',
		WEB=>'0',
		SSRB=>'0',
		ADDRB=>AD2(10 downto 0),
		DIB=>(others=>'0'),
		DIPB(0)=>'0',
		DOB=>doutb(2)(15 downto 8),
		DOPB(0)=>pout(11)
	);
	
	XLXI_6 : RAMB16_S9_S9
	generic map (
		INIT_00=>cRAMDoublePort_XLXI_6_INIT_00,
		INIT_01=>cRAMDoublePort_XLXI_6_INIT_01,
		INIT_02=>cRAMDoublePort_XLXI_6_INIT_02,
		INIT_03=>cRAMDoublePort_XLXI_6_INIT_03,
		INIT_04=>cRAMDoublePort_XLXI_6_INIT_04,
		INIT_05=>cRAMDoublePort_XLXI_6_INIT_05,
		INIT_06=>cRAMDoublePort_XLXI_6_INIT_06,
		INIT_07=>cRAMDoublePort_XLXI_6_INIT_07,
		INIT_08=>cRAMDoublePort_XLXI_6_INIT_08,
		INIT_09=>cRAMDoublePort_XLXI_6_INIT_09,
		INIT_0a=>cRAMDoublePort_XLXI_6_INIT_0A,
		INIT_0b=>cRAMDoublePort_XLXI_6_INIT_0B,
		INIT_0c=>cRAMDoublePort_XLXI_6_INIT_0C,
		INIT_0d=>cRAMDoublePort_XLXI_6_INIT_0D,
		INIT_0e=>cRAMDoublePort_XLXI_6_INIT_0E,
		INIT_0f=>cRAMDoublePort_XLXI_6_INIT_0F,
		INIT_10=>cRAMDoublePort_XLXI_6_INIT_10,
		INIT_11=>cRAMDoublePort_XLXI_6_INIT_11,
		INIT_12=>cRAMDoublePort_XLXI_6_INIT_12,
		INIT_13=>cRAMDoublePort_XLXI_6_INIT_13,
		INIT_14=>cRAMDoublePort_XLXI_6_INIT_14,
		INIT_15=>cRAMDoublePort_XLXI_6_INIT_15,
		INIT_16=>cRAMDoublePort_XLXI_6_INIT_16,
		INIT_17=>cRAMDoublePort_XLXI_6_INIT_17,
		INIT_18=>cRAMDoublePort_XLXI_6_INIT_18,
		INIT_19=>cRAMDoublePort_XLXI_6_INIT_19,
		INIT_1a=>cRAMDoublePort_XLXI_6_INIT_1A,
		INIT_1b=>cRAMDoublePort_XLXI_6_INIT_1B,
		INIT_1c=>cRAMDoublePort_XLXI_6_INIT_1C,
		INIT_1d=>cRAMDoublePort_XLXI_6_INIT_1D,
		INIT_1e=>cRAMDoublePort_XLXI_6_INIT_1E,
		INIT_1f=>cRAMDoublePort_XLXI_6_INIT_1F,
		INIT_20=>cRAMDoublePort_XLXI_6_INIT_20,
		INIT_21=>cRAMDoublePort_XLXI_6_INIT_21,
		INIT_22=>cRAMDoublePort_XLXI_6_INIT_22,
		INIT_23=>cRAMDoublePort_XLXI_6_INIT_23,
		INIT_24=>cRAMDoublePort_XLXI_6_INIT_24,
		INIT_25=>cRAMDoublePort_XLXI_6_INIT_25,
		INIT_26=>cRAMDoublePort_XLXI_6_INIT_26,
		INIT_27=>cRAMDoublePort_XLXI_6_INIT_27,
		INIT_28=>cRAMDoublePort_XLXI_6_INIT_28,
		INIT_29=>cRAMDoublePort_XLXI_6_INIT_29,
		INIT_2a=>cRAMDoublePort_XLXI_6_INIT_2A,
		INIT_2b=>cRAMDoublePort_XLXI_6_INIT_2B,
		INIT_2c=>cRAMDoublePort_XLXI_6_INIT_2C,
		INIT_2d=>cRAMDoublePort_XLXI_6_INIT_2D,
		INIT_2e=>cRAMDoublePort_XLXI_6_INIT_2E,
		INIT_2f=>cRAMDoublePort_XLXI_6_INIT_2F,
		INIT_30=>cRAMDoublePort_XLXI_6_INIT_30,
		INIT_31=>cRAMDoublePort_XLXI_6_INIT_31,
		INIT_32=>cRAMDoublePort_XLXI_6_INIT_32,
		INIT_33=>cRAMDoublePort_XLXI_6_INIT_33,
		INIT_34=>cRAMDoublePort_XLXI_6_INIT_34,
		INIT_35=>cRAMDoublePort_XLXI_6_INIT_35,
		INIT_36=>cRAMDoublePort_XLXI_6_INIT_36,
		INIT_37=>cRAMDoublePort_XLXI_6_INIT_37,
		INIT_38=>cRAMDoublePort_XLXI_6_INIT_38,
		INIT_39=>cRAMDoublePort_XLXI_6_INIT_39,
		INIT_3a=>cRAMDoublePort_XLXI_6_INIT_3A,
		INIT_3b=>cRAMDoublePort_XLXI_6_INIT_3B,
		INIT_3c=>cRAMDoublePort_XLXI_6_INIT_3C,
		INIT_3d=>cRAMDoublePort_XLXI_6_INIT_3D,
		INIT_3e=>cRAMDoublePort_XLXI_6_INIT_3E,
		INIT_3f=>cRAMDoublePort_XLXI_6_INIT_3F
	)
	port map (
		CLKA=>CLK,
		ENA=>CE1,
		WEA=>WE1,
		SSRA=>'0',
		ADDRA=>AD1(10 downto 0),
		DIA=>DIN1(7 downto 0),
		DIPA(0)=>plow,
		DOA=>douta(3)(7 downto 0),
		DOPA(0)=>pout(12),
		
		CLKB=>CLK,
		ENB=>'1',
		WEB=>'0',
		SSRB=>'0',
		ADDRB=>AD2(10 downto 0),
		DIB=>(others=>'0'),
		DIPB(0)=>'0',
		DOB=>doutb(3)(7 downto 0),
		DOPB(0)=>pout(13)
	);
	
	XLXI_7 : RAMB16_S9_S9
	generic map (
		INIT_00=>cRAMDoublePort_XLXI_7_INIT_00,
		INIT_01=>cRAMDoublePort_XLXI_7_INIT_01,
		INIT_02=>cRAMDoublePort_XLXI_7_INIT_02,
		INIT_03=>cRAMDoublePort_XLXI_7_INIT_03,
		INIT_04=>cRAMDoublePort_XLXI_7_INIT_04,
		INIT_05=>cRAMDoublePort_XLXI_7_INIT_05,
		INIT_06=>cRAMDoublePort_XLXI_7_INIT_06,
		INIT_07=>cRAMDoublePort_XLXI_7_INIT_07,
		INIT_08=>cRAMDoublePort_XLXI_7_INIT_08,
		INIT_09=>cRAMDoublePort_XLXI_7_INIT_09,
		INIT_0a=>cRAMDoublePort_XLXI_7_INIT_0A,
		INIT_0b=>cRAMDoublePort_XLXI_7_INIT_0B,
		INIT_0c=>cRAMDoublePort_XLXI_7_INIT_0C,
		INIT_0d=>cRAMDoublePort_XLXI_7_INIT_0D,
		INIT_0e=>cRAMDoublePort_XLXI_7_INIT_0E,
		INIT_0f=>cRAMDoublePort_XLXI_7_INIT_0F,
		INIT_10=>cRAMDoublePort_XLXI_7_INIT_10,
		INIT_11=>cRAMDoublePort_XLXI_7_INIT_11,
		INIT_12=>cRAMDoublePort_XLXI_7_INIT_12,
		INIT_13=>cRAMDoublePort_XLXI_7_INIT_13,
		INIT_14=>cRAMDoublePort_XLXI_7_INIT_14,
		INIT_15=>cRAMDoublePort_XLXI_7_INIT_15,
		INIT_16=>cRAMDoublePort_XLXI_7_INIT_16,
		INIT_17=>cRAMDoublePort_XLXI_7_INIT_17,
		INIT_18=>cRAMDoublePort_XLXI_7_INIT_18,
		INIT_19=>cRAMDoublePort_XLXI_7_INIT_19,
		INIT_1a=>cRAMDoublePort_XLXI_7_INIT_1A,
		INIT_1b=>cRAMDoublePort_XLXI_7_INIT_1B,
		INIT_1c=>cRAMDoublePort_XLXI_7_INIT_1C,
		INIT_1d=>cRAMDoublePort_XLXI_7_INIT_1D,
		INIT_1e=>cRAMDoublePort_XLXI_7_INIT_1E,
		INIT_1f=>cRAMDoublePort_XLXI_7_INIT_1F,
		INIT_20=>cRAMDoublePort_XLXI_7_INIT_20,
		INIT_21=>cRAMDoublePort_XLXI_7_INIT_21,
		INIT_22=>cRAMDoublePort_XLXI_7_INIT_22,
		INIT_23=>cRAMDoublePort_XLXI_7_INIT_23,
		INIT_24=>cRAMDoublePort_XLXI_7_INIT_24,
		INIT_25=>cRAMDoublePort_XLXI_7_INIT_25,
		INIT_26=>cRAMDoublePort_XLXI_7_INIT_26,
		INIT_27=>cRAMDoublePort_XLXI_7_INIT_27,
		INIT_28=>cRAMDoublePort_XLXI_7_INIT_28,
		INIT_29=>cRAMDoublePort_XLXI_7_INIT_29,
		INIT_2a=>cRAMDoublePort_XLXI_7_INIT_2A,
		INIT_2b=>cRAMDoublePort_XLXI_7_INIT_2B,
		INIT_2c=>cRAMDoublePort_XLXI_7_INIT_2C,
		INIT_2d=>cRAMDoublePort_XLXI_7_INIT_2D,
		INIT_2e=>cRAMDoublePort_XLXI_7_INIT_2E,
		INIT_2f=>cRAMDoublePort_XLXI_7_INIT_2F,
		INIT_30=>cRAMDoublePort_XLXI_7_INIT_30,
		INIT_31=>cRAMDoublePort_XLXI_7_INIT_31,
		INIT_32=>cRAMDoublePort_XLXI_7_INIT_32,
		INIT_33=>cRAMDoublePort_XLXI_7_INIT_33,
		INIT_34=>cRAMDoublePort_XLXI_7_INIT_34,
		INIT_35=>cRAMDoublePort_XLXI_7_INIT_35,
		INIT_36=>cRAMDoublePort_XLXI_7_INIT_36,
		INIT_37=>cRAMDoublePort_XLXI_7_INIT_37,
		INIT_38=>cRAMDoublePort_XLXI_7_INIT_38,
		INIT_39=>cRAMDoublePort_XLXI_7_INIT_39,
		INIT_3a=>cRAMDoublePort_XLXI_7_INIT_3A,
		INIT_3b=>cRAMDoublePort_XLXI_7_INIT_3B,
		INIT_3c=>cRAMDoublePort_XLXI_7_INIT_3C,
		INIT_3d=>cRAMDoublePort_XLXI_7_INIT_3D,
		INIT_3e=>cRAMDoublePort_XLXI_7_INIT_3E,
		INIT_3f=>cRAMDoublePort_XLXI_7_INIT_3F
	)
	port map (
		CLKA=>CLK,
		ENA=>CE1,
		WEA=>WE1,
		SSRA=>'0',
		ADDRA=>AD1(10 downto 0),
		DIA=>DIN1(15 downto 8),
		DIPA(0)=>phigh,
		DOA=>douta(3)(15 downto 8),
		DOPA(0)=>pout(14),
		
		CLKB=>CLK,
		ENB=>'1',
		WEB=>'0',
		SSRB=>'0',
		ADDRB=>AD2(10 downto 0),
		DIB=>(others=>'0'),
		DIPB(0)=>'0',
		DOB=>doutb(3)(15 downto 8),
		DOPB(0)=>pout(15)
	);
	
	DOUT1 <= douta(to_integer(unsigned(AD1(12 downto 11))));
	DOUT2 <= doutb(to_integer(unsigned(AD2(12 downto 11))));
end BEHAVIORAL;
