----------------------------------------------------------------------------------
--
-- File retrieved, on 07/02/2010, from :
-- http://sebastien-viardot.imag.fr/Enseignements/Archi1A2s/sources/RAMDoublePort.vhd
--
-- Slightly altered to get rid of vendor-specific packages and adjust formatting
--
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity RAMDoublePort is
    Port ( AD1 : in  STD_LOGIC_VECTOR (12 downto 0);
           AD2 : in  STD_LOGIC_VECTOR (12 downto 0);
           DIN1 : in  STD_LOGIC_VECTOR (15 downto 0);
           DOUT1 : out  STD_LOGIC_VECTOR (15 downto 0);
           WE1 : in  STD_LOGIC;
           DOUT2 : out  STD_LOGIC_VECTOR (15 downto 0);
           OE1 : in  STD_LOGIC;
           CE1 : in  STD_LOGIC;
			  CLK : in STD_LOGIC);
end RAMDoublePort;

 -- memory map :
 --     0 -  4799 : VGA-mapped RAM (320*240 pix, 16 pix per word => 4800 words)
 --  4800 -  5823 : font map (8*8 : 4 words per character, 256 chars => 1024 words)
 --  5824 -  8191 : user data (2368 words)

architecture Behavioral of RAMDoublePort is
 constant low_address: natural := 0;
 constant high_address: natural := 8192;  
 subtype octet is std_logic_vector( 15 downto 0 );
 type zone_memoire is
         array (natural range low_address to high_address) of octet;
 signal memoire: zone_memoire := (
 -- 0 - 4799 : VGA-mapped RAM
 
 -- 4800 - 5823  : font map (8*8 : 4 words per character, 256 chars => 1024 words)
   4800=> "00000000"
        & "00000000",
   4801=> "00000000"
        & "00000000",
   4802=> "00000000"
        & "00000000",
   4803=> "00000000"
        & "00000000",
   4804=> "00000000"
        & "01010000",
   4805=> "00000000"
        & "00000000",
   4806=> "10001000"
        & "01110000",
   4807=> "00000000"
        & "00000000",
   4808=> "00000000"
        & "01010000",
   4809=> "00000000"
        & "00000000",
   4810=> "01110000"
        & "10001000",
   4811=> "00000000"
        & "00000000",
   4812=> "01010000"
        & "11111000",
   4813=> "11111000"
        & "11111000",
   4814=> "11111000"
        & "01110000",
   4815=> "00100000"
        & "00000000",
   4816=> "00100000"
        & "01110000",
   4817=> "11111000"
        & "11111000",
   4818=> "11111000"
        & "01110000",
   4819=> "00100000"
        & "00000000",
   4820=> "01110000"
        & "01110000",
   4821=> "00100000"
        & "11111000",
   4822=> "11111000"
        & "00100000",
   4823=> "01110000"
        & "00000000",
   4824=> "00100000"
        & "01110000",
   4825=> "11111000"
        & "11111000",
   4826=> "01110000"
        & "00100000",
   4827=> "01110000"
        & "00000000",
   4828=> "00000000"
        & "00000000",
   4829=> "01110000"
        & "01110000",
   4830=> "01110000"
        & "00000000",
   4831=> "00000000"
        & "00000000",
   4832=> "11111000"
        & "11111000",
   4833=> "10001000"
        & "10001000",
   4834=> "10001000"
        & "11111000",
   4835=> "11111000"
        & "00000000",
   4836=> "00000000"
        & "00000000",
   4837=> "01110000"
        & "01010000",
   4838=> "01110000"
        & "00000000",
   4839=> "00000000"
        & "00000000",
   4840=> "11111000"
        & "11111000",
   4841=> "10001000"
        & "10101000",
   4842=> "10001000"
        & "11111000",
   4843=> "11111000"
        & "00000000",
   4844=> "00100000"
        & "01110000",
   4845=> "10101000"
        & "00100000",
   4846=> "01110000"
        & "10001000",
   4847=> "01110000"
        & "00000000",
   4848=> "01110000"
        & "10001000",
   4849=> "01110000"
        & "00100000",
   4850=> "00100000"
        & "11111000",
   4851=> "00100000"
        & "00000000",
   4852=> "00111000"
        & "00111000",
   4853=> "00100000"
        & "00100000",
   4854=> "01100000"
        & "11100000",
   4855=> "01100000"
        & "00000000",
   4856=> "01111000"
        & "01111000",
   4857=> "01001000"
        & "01011000",
   4858=> "01011000"
        & "11000000",
   4859=> "11000000"
        & "00000000",
   4860=> "00000000"
        & "10101000",
   4861=> "01010000"
        & "10001000",
   4862=> "01010000"
        & "10101000",
   4863=> "00000000"
        & "00000000",
   4864=> "01000000"
        & "01100000",
   4865=> "01110000"
        & "01111000",
   4866=> "01110000"
        & "01100000",
   4867=> "01000000"
        & "00000000",
   4868=> "00010000"
        & "00110000",
   4869=> "01110000"
        & "11110000",
   4870=> "01110000"
        & "00110000",
   4871=> "00010000"
        & "00000000",
   4872=> "00100000"
        & "01110000",
   4873=> "10101000"
        & "00100000",
   4874=> "10101000"
        & "01110000",
   4875=> "00100000"
        & "00000000",
   4876=> "01010000"
        & "01010000",
   4877=> "01010000"
        & "01010000",
   4878=> "00000000"
        & "01010000",
   4879=> "01010000"
        & "00000000",
   4880=> "01111000"
        & "11101000",
   4881=> "11101000"
        & "01111000",
   4882=> "00101000"
        & "00101000",
   4883=> "00101000"
        & "00000000",
   4884=> "01111000"
        & "11001000",
   4885=> "10100000"
        & "01010000",
   4886=> "00101000"
        & "10011000",
   4887=> "11110000"
        & "00000000",
   4888=> "00000000"
        & "00000000",
   4889=> "00000000"
        & "00000000",
   4890=> "11111000"
        & "11111000",
   4891=> "11111000"
        & "00000000",
   4892=> "00100000"
        & "01110000",
   4893=> "00100000"
        & "00100000",
   4894=> "01110000"
        & "00100000",
   4895=> "11111000"
        & "00000000",
   4896=> "00100000"
        & "01110000",
   4897=> "11111000"
        & "00100000",
   4898=> "00100000"
        & "00100000",
   4899=> "00100000"
        & "00000000",
   4900=> "00100000"
        & "00100000",
   4901=> "00100000"
        & "00100000",
   4902=> "11111000"
        & "01110000",
   4903=> "00100000"
        & "00000000",
   4904=> "00000000"
        & "00100000",
   4905=> "00110000"
        & "11111000",
   4906=> "00110000"
        & "00100000",
   4907=> "00000000"
        & "00000000",
   4908=> "00000000"
        & "00100000",
   4909=> "01100000"
        & "11111000",
   4910=> "01100000"
        & "00100000",
   4911=> "00000000"
        & "00000000",
   4912=> "00000000"
        & "00000000",
   4913=> "01000000"
        & "01111000",
   4914=> "00000000"
        & "00000000",
   4915=> "00000000"
        & "00000000",
   4916=> "00000000"
        & "00000000",
   4917=> "01010000"
        & "11111000",
   4918=> "01010000"
        & "00000000",
   4919=> "00000000"
        & "00000000",
   4920=> "00000000"
        & "00100000",
   4921=> "00100000"
        & "01110000",
   4922=> "01110000"
        & "11111000",
   4923=> "11111000"
        & "00000000",
   4924=> "11111000"
        & "11111000",
   4925=> "01110000"
        & "01110000",
   4926=> "00100000"
        & "00100000",
   4927=> "00000000"
        & "00000000",
   4928=> "00000000"
        & "00000000",
   4929=> "00000000"
        & "00000000",
   4930=> "00000000"
        & "00000000",
   4931=> "00000000"
        & "00000000",
   4932=> "00100000"
        & "00100000",
   4933=> "00100000"
        & "00100000",
   4934=> "00000000"
        & "00100000",
   4935=> "00100000"
        & "00000000",
   4936=> "01010000"
        & "01010000",
   4937=> "01010000"
        & "00000000",
   4938=> "00000000"
        & "00000000",
   4939=> "00000000"
        & "00000000",
   4940=> "01010000"
        & "01010000",
   4941=> "11111000"
        & "01010000",
   4942=> "11111000"
        & "01010000",
   4943=> "01010000"
        & "00000000",
   4944=> "00100000"
        & "01110000",
   4945=> "10100000"
        & "01110000",
   4946=> "00101000"
        & "01110000",
   4947=> "00100000"
        & "00000000",
   4948=> "11000000"
        & "11001000",
   4949=> "00010000"
        & "00100000",
   4950=> "01000000"
        & "10011000",
   4951=> "00011000"
        & "00000000",
   4952=> "01000000"
        & "10100000",
   4953=> "10100000"
        & "01000000",
   4954=> "10101000"
        & "10010000",
   4955=> "01101000"
        & "00000000",
   4956=> "00100000"
        & "00100000",
   4957=> "01000000"
        & "00000000",
   4958=> "00000000"
        & "00000000",
   4959=> "00000000"
        & "00000000",
   4960=> "00010000"
        & "00100000",
   4961=> "01000000"
        & "01000000",
   4962=> "01000000"
        & "00100000",
   4963=> "00010000"
        & "00000000",
   4964=> "01000000"
        & "00100000",
   4965=> "00010000"
        & "00010000",
   4966=> "00010000"
        & "00100000",
   4967=> "01000000"
        & "00000000",
   4968=> "10101000"
        & "01110000",
   4969=> "10101000"
        & "00000000",
   4970=> "00000000"
        & "00000000",
   4971=> "00000000"
        & "00000000",
   4972=> "00000000"
        & "00100000",
   4973=> "00100000"
        & "11111000",
   4974=> "00100000"
        & "00100000",
   4975=> "00000000"
        & "00000000",
   4976=> "00000000"
        & "00000000",
   4977=> "00000000"
        & "00000000",
   4978=> "01100000"
        & "00100000",
   4979=> "01000000"
        & "00000000",
   4980=> "00000000"
        & "00000000",
   4981=> "00000000"
        & "11111000",
   4982=> "00000000"
        & "00000000",
   4983=> "00000000"
        & "00000000",
   4984=> "00000000"
        & "00000000",
   4985=> "00000000"
        & "00000000",
   4986=> "00000000"
        & "01100000",
   4987=> "01100000"
        & "00000000",
   4988=> "00000000"
        & "00001000",
   4989=> "00010000"
        & "00100000",
   4990=> "01000000"
        & "10000000",
   4991=> "00000000"
        & "00000000",
   4992=> "01110000"
        & "10001000",
   4993=> "10011000"
        & "10101000",
   4994=> "11001000"
        & "10001000",
   4995=> "01110000"
        & "00000000",
   4996=> "00100000"
        & "11100000",
   4997=> "00100000"
        & "00100000",
   4998=> "00100000"
        & "00100000",
   4999=> "11111000"
        & "00000000",
   5000=> "01110000"
        & "10001000",
   5001=> "00001000"
        & "00110000",
   5002=> "01000000"
        & "10000000",
   5003=> "11111000"
        & "00000000",
   5004=> "01110000"
        & "10001000",
   5005=> "00001000"
        & "00110000",
   5006=> "00001000"
        & "10001000",
   5007=> "01110000"
        & "00000000",
   5008=> "10001000"
        & "10001000",
   5009=> "10001000"
        & "11111000",
   5010=> "00001000"
        & "00001000",
   5011=> "00001000"
        & "00000000",
   5012=> "11111000"
        & "10000000",
   5013=> "11110000"
        & "00001000",
   5014=> "00001000"
        & "10001000",
   5015=> "01110000"
        & "00000000",
   5016=> "01110000"
        & "10000000",
   5017=> "10000000"
        & "11110000",
   5018=> "10001000"
        & "10001000",
   5019=> "01110000"
        & "00000000",
   5020=> "11111000"
        & "00001000",
   5021=> "00001000"
        & "00010000",
   5022=> "00100000"
        & "00100000",
   5023=> "00100000"
        & "00000000",
   5024=> "01110000"
        & "10001000",
   5025=> "10001000"
        & "01110000",
   5026=> "10001000"
        & "10001000",
   5027=> "01110000"
        & "00000000",
   5028=> "01110000"
        & "10001000",
   5029=> "10001000"
        & "01111000",
   5030=> "00001000"
        & "00001000",
   5031=> "01110000"
        & "00000000",
   5032=> "00000000"
        & "01100000",
   5033=> "01100000"
        & "00000000",
   5034=> "01100000"
        & "01100000",
   5035=> "00000000"
        & "00000000",
   5036=> "00000000"
        & "01100000",
   5037=> "01100000"
        & "00000000",
   5038=> "01100000"
        & "00100000",
   5039=> "01000000"
        & "00000000",
   5040=> "00010000"
        & "00100000",
   5041=> "01000000"
        & "10000000",
   5042=> "01000000"
        & "00100000",
   5043=> "00010000"
        & "00000000",
   5044=> "00000000"
        & "00000000",
   5045=> "11111000"
        & "00000000",
   5046=> "11111000"
        & "00000000",
   5047=> "00000000"
        & "00000000",
   5048=> "01000000"
        & "00100000",
   5049=> "00010000"
        & "00001000",
   5050=> "00010000"
        & "00100000",
   5051=> "01000000"
        & "00000000",
   5052=> "01110000"
        & "10001000",
   5053=> "00001000"
        & "00010000",
   5054=> "00100000"
        & "00000000",
   5055=> "00100000"
        & "00000000",
   5056=> "01110000"
        & "10001000",
   5057=> "10011000"
        & "10101000",
   5058=> "10011000"
        & "10000000",
   5059=> "01110000"
        & "00000000",
   5060=> "00100000"
        & "00100000",
   5061=> "01010000"
        & "01110000",
   5062=> "01010000"
        & "10001000",
   5063=> "10001000"
        & "00000000",
   5064=> "11110000"
        & "10001000",
   5065=> "10001000"
        & "11110000",
   5066=> "10001000"
        & "10001000",
   5067=> "11110000"
        & "00000000",
   5068=> "01110000"
        & "10001000",
   5069=> "10000000"
        & "10000000",
   5070=> "10000000"
        & "10001000",
   5071=> "01110000"
        & "00000000",
   5072=> "11110000"
        & "10001000",
   5073=> "10001000"
        & "10001000",
   5074=> "10001000"
        & "10001000",
   5075=> "11110000"
        & "00000000",
   5076=> "11111000"
        & "10000000",
   5077=> "10000000"
        & "11110000",
   5078=> "10000000"
        & "10000000",
   5079=> "11111000"
        & "00000000",
   5080=> "11111000"
        & "10000000",
   5081=> "10000000"
        & "11110000",
   5082=> "10000000"
        & "10000000",
   5083=> "10000000"
        & "00000000",
   5084=> "01110000"
        & "10001000",
   5085=> "10000000"
        & "10111000",
   5086=> "10001000"
        & "10001000",
   5087=> "01110000"
        & "00000000",
   5088=> "10001000"
        & "10001000",
   5089=> "10001000"
        & "11111000",
   5090=> "10001000"
        & "10001000",
   5091=> "10001000"
        & "00000000",
   5092=> "11111000"
        & "00100000",
   5093=> "00100000"
        & "00100000",
   5094=> "00100000"
        & "00100000",
   5095=> "11111000"
        & "00000000",
   5096=> "00001000"
        & "00001000",
   5097=> "00001000"
        & "00001000",
   5098=> "00001000"
        & "10001000",
   5099=> "01110000"
        & "00000000",
   5100=> "10001000"
        & "10010000",
   5101=> "10100000"
        & "11000000",
   5102=> "10100000"
        & "10010000",
   5103=> "10001000"
        & "00000000",
   5104=> "10000000"
        & "10000000",
   5105=> "10000000"
        & "10000000",
   5106=> "10000000"
        & "10000000",
   5107=> "11111000"
        & "00000000",
   5108=> "10001000"
        & "11011000",
   5109=> "10101000"
        & "10001000",
   5110=> "10001000"
        & "10001000",
   5111=> "10001000"
        & "00000000",
   5112=> "10001000"
        & "11001000",
   5113=> "10101000"
        & "10011000",
   5114=> "10001000"
        & "10001000",
   5115=> "10001000"
        & "00000000",
   5116=> "01110000"
        & "10001000",
   5117=> "10001000"
        & "10001000",
   5118=> "10001000"
        & "10001000",
   5119=> "01110000"
        & "00000000",
   5120=> "11110000"
        & "10001000",
   5121=> "10001000"
        & "11110000",
   5122=> "10000000"
        & "10000000",
   5123=> "10000000"
        & "00000000",
   5124=> "01110000"
        & "10001000",
   5125=> "10001000"
        & "10001000",
   5126=> "10101000"
        & "10010000",
   5127=> "01101000"
        & "00000000",
   5128=> "11110000"
        & "10001000",
   5129=> "10001000"
        & "11110000",
   5130=> "10010000"
        & "10001000",
   5131=> "10001000"
        & "00000000",
   5132=> "01110000"
        & "10001000",
   5133=> "10000000"
        & "01110000",
   5134=> "00001000"
        & "10001000",
   5135=> "01110000"
        & "00000000",
   5136=> "11111000"
        & "00100000",
   5137=> "00100000"
        & "00100000",
   5138=> "00100000"
        & "00100000",
   5139=> "00100000"
        & "00000000",
   5140=> "10001000"
        & "10001000",
   5141=> "10001000"
        & "10001000",
   5142=> "10001000"
        & "10001000",
   5143=> "01110000"
        & "00000000",
   5144=> "10001000"
        & "10001000",
   5145=> "10001000"
        & "10001000",
   5146=> "10001000"
        & "01010000",
   5147=> "00100000"
        & "00000000",
   5148=> "10001000"
        & "10001000",
   5149=> "10001000"
        & "10001000",
   5150=> "10101000"
        & "11011000",
   5151=> "10001000"
        & "00000000",
   5152=> "10001000"
        & "10001000",
   5153=> "01010000"
        & "00100000",
   5154=> "01010000"
        & "10001000",
   5155=> "10001000"
        & "00000000",
   5156=> "10001000"
        & "10001000",
   5157=> "10001000"
        & "01010000",
   5158=> "00100000"
        & "00100000",
   5159=> "00100000"
        & "00000000",
   5160=> "11111000"
        & "00001000",
   5161=> "00010000"
        & "00100000",
   5162=> "01000000"
        & "10000000",
   5163=> "11111000"
        & "00000000",
   5164=> "01110000"
        & "01000000",
   5165=> "01000000"
        & "01000000",
   5166=> "01000000"
        & "01000000",
   5167=> "01110000"
        & "00000000",
   5168=> "00000000"
        & "10000000",
   5169=> "01000000"
        & "00100000",
   5170=> "00010000"
        & "00001000",
   5171=> "00000000"
        & "00000000",
   5172=> "01110000"
        & "00010000",
   5173=> "00010000"
        & "00010000",
   5174=> "00010000"
        & "00010000",
   5175=> "01110000"
        & "00000000",
   5176=> "00100000"
        & "01010000",
   5177=> "10001000"
        & "00000000",
   5178=> "00000000"
        & "00000000",
   5179=> "00000000"
        & "00000000",
   5180=> "00000000"
        & "00000000",
   5181=> "00000000"
        & "00000000",
   5182=> "00000000"
        & "00000000",
   5183=> "11111000"
        & "00000000",
   5184=> "00000000"
        & "00010000",
   5185=> "00100000"
        & "00000000",
   5186=> "00000000"
        & "00000000",
   5187=> "00000000"
        & "00000000",
   5188=> "00000000"
        & "00000000",
   5189=> "01110000"
        & "00001000",
   5190=> "01111000"
        & "10001000",
   5191=> "01111000"
        & "00000000",
   5192=> "10000000"
        & "10000000",
   5193=> "10000000"
        & "11110000",
   5194=> "10001000"
        & "10001000",
   5195=> "11110000"
        & "00000000",
   5196=> "00000000"
        & "00000000",
   5197=> "01110000"
        & "10001000",
   5198=> "10000000"
        & "10001000",
   5199=> "01110000"
        & "00000000",
   5200=> "00001000"
        & "00001000",
   5201=> "00001000"
        & "01111000",
   5202=> "10001000"
        & "10001000",
   5203=> "01111000"
        & "00000000",
   5204=> "00000000"
        & "00000000",
   5205=> "01110000"
        & "10001000",
   5206=> "11111000"
        & "10000000",
   5207=> "01111000"
        & "00000000",
   5208=> "00110000"
        & "01001000",
   5209=> "01000000"
        & "11100000",
   5210=> "01000000"
        & "01000000",
   5211=> "01000000"
        & "00000000",
   5212=> "00000000"
        & "00000000",
   5213=> "01111000"
        & "10001000",
   5214=> "01111000"
        & "00001000",
   5215=> "11110000"
        & "00000000",
   5216=> "10000000"
        & "10000000",
   5217=> "10000000"
        & "11110000",
   5218=> "10001000"
        & "10001000",
   5219=> "10001000"
        & "00000000",
   5220=> "00000000"
        & "00100000",
   5221=> "00000000"
        & "01100000",
   5222=> "00100000"
        & "00100000",
   5223=> "01110000"
        & "00000000",
   5224=> "00000000"
        & "00010000",
   5225=> "00000000"
        & "00010000",
   5226=> "00010000"
        & "10010000",
   5227=> "01100000"
        & "00000000",
   5228=> "10000000"
        & "10000000",
   5229=> "10010000"
        & "10100000",
   5230=> "11000000"
        & "10100000",
   5231=> "10011000"
        & "00000000",
   5232=> "01100000"
        & "00100000",
   5233=> "00100000"
        & "00100000",
   5234=> "00100000"
        & "00100000",
   5235=> "01110000"
        & "00000000",
   5236=> "00000000"
        & "00000000",
   5237=> "11010000"
        & "10101000",
   5238=> "10101000"
        & "10001000",
   5239=> "10001000"
        & "00000000",
   5240=> "00000000"
        & "00000000",
   5241=> "10110000"
        & "11001000",
   5242=> "10001000"
        & "10001000",
   5243=> "10001000"
        & "00000000",
   5244=> "00000000"
        & "00000000",
   5245=> "01110000"
        & "10001000",
   5246=> "10001000"
        & "10001000",
   5247=> "01110000"
        & "00000000",
   5248=> "00000000"
        & "00000000",
   5249=> "11110000"
        & "10001000",
   5250=> "11110000"
        & "10000000",
   5251=> "10000000"
        & "00000000",
   5252=> "00000000"
        & "00000000",
   5253=> "01111000"
        & "10001000",
   5254=> "01111000"
        & "00001000",
   5255=> "00001000"
        & "00000000",
   5256=> "00000000"
        & "00000000",
   5257=> "10110000"
        & "11001000",
   5258=> "10000000"
        & "10000000",
   5259=> "10000000"
        & "00000000",
   5260=> "00000000"
        & "00000000",
   5261=> "01111000"
        & "10000000",
   5262=> "01110000"
        & "00001000",
   5263=> "11110000"
        & "00000000",
   5264=> "01000000"
        & "01000000",
   5265=> "11100000"
        & "01000000",
   5266=> "01000000"
        & "01001000",
   5267=> "00110000"
        & "00000000",
   5268=> "00000000"
        & "00000000",
   5269=> "10001000"
        & "10001000",
   5270=> "10001000"
        & "10011000",
   5271=> "01101000"
        & "00000000",
   5272=> "00000000"
        & "00000000",
   5273=> "10001000"
        & "10001000",
   5274=> "10001000"
        & "01010000",
   5275=> "00100000"
        & "00000000",
   5276=> "00000000"
        & "00000000",
   5277=> "10001000"
        & "10001000",
   5278=> "10001000"
        & "10101000",
   5279=> "01010000"
        & "00000000",
   5280=> "00000000"
        & "00000000",
   5281=> "10001000"
        & "01010000",
   5282=> "00100000"
        & "01010000",
   5283=> "10001000"
        & "00000000",
   5284=> "00000000"
        & "00000000",
   5285=> "10001000"
        & "01010000",
   5286=> "00100000"
        & "01000000",
   5287=> "10000000"
        & "00000000",
   5288=> "00000000"
        & "00000000",
   5289=> "11111000"
        & "00010000",
   5290=> "00100000"
        & "01000000",
   5291=> "11111000"
        & "00000000",
   5292=> "00011000"
        & "00100000",
   5293=> "00100000"
        & "01000000",
   5294=> "00100000"
        & "00100000",
   5295=> "00011000"
        & "00000000",
   5296=> "00100000"
        & "00100000",
   5297=> "00100000"
        & "00000000",
   5298=> "00100000"
        & "00100000",
   5299=> "00100000"
        & "00000000",
   5300=> "01100000"
        & "00010000",
   5301=> "00010000"
        & "00001000",
   5302=> "00010000"
        & "00010000",
   5303=> "01100000"
        & "00000000",
   5304=> "00000000"
        & "00000000",
   5305=> "01000000"
        & "10101000",
   5306=> "00010000"
        & "00000000",
   5307=> "00000000"
        & "00000000",
   5308=> "00000000"
        & "00100000",
   5309=> "01010000"
        & "10001000",
   5310=> "10001000"
        & "10001000",
   5311=> "11111000"
        & "00000000",
   5312=> "01110000"
        & "10001000",
   5313=> "10000000"
        & "10001000",
   5314=> "01110000"
        & "00100000",
   5315=> "11000000"
        & "00000000",
   5316=> "00000000"
        & "01110000",
   5317=> "10000000"
        & "10001000",
   5318=> "01110000"
        & "00100000",
   5319=> "11000000"
        & "00000000",
   5320=> "00010100"
        & "01001000",
   5321=> "10001000"
        & "11001000",
   5322=> "10101000"
        & "10011000",
   5323=> "10001000"
        & "00000000",
   5324=> "00101000"
        & "01010000",
   5325=> "00000000"
        & "10110000",
   5326=> "11001000"
        & "10001000",
   5327=> "10001000"
        & "00000000",
   5328=> "00010000"
        & "00100000",
   5329=> "01110000"
        & "10001000",
   5330=> "11111000"
        & "10001000",
   5331=> "10001000"
        & "00000000",
   5332=> "01000000"
        & "00100000",
   5333=> "01110000"
        & "10001000",
   5334=> "11111000"
        & "10001000",
   5335=> "10001000"
        & "00000000",
   5336=> "01010000"
        & "00000000",
   5337=> "01110000"
        & "10001000",
   5338=> "11111000"
        & "10001000",
   5339=> "10001000"
        & "00000000",
   5340=> "00100000"
        & "01010000",
   5341=> "00000000"
        & "01110000",
   5342=> "10001000"
        & "11111000",
   5343=> "10001000"
        & "00000000",
   5344=> "00010000"
        & "00100000",
   5345=> "11111000"
        & "10000000",
   5346=> "11110000"
        & "10000000",
   5347=> "11111000"
        & "00000000",
   5348=> "01000000"
        & "00100000",
   5349=> "11111000"
        & "10000000",
   5350=> "11110000"
        & "10000000",
   5351=> "11111000"
        & "00000000",
   5352=> "01010000"
        & "00000000",
   5353=> "11111000"
        & "10000000",
   5354=> "11110000"
        & "10000000",
   5355=> "11111000"
        & "00000000",
   5356=> "00100000"
        & "01010000",
   5357=> "11111000"
        & "10000000",
   5358=> "11110000"
        & "10000000",
   5359=> "11111000"
        & "00000000",
   5360=> "00010000"
        & "00100000",
   5361=> "11111000"
        & "00100000",
   5362=> "00100000"
        & "00100000",
   5363=> "11111000"
        & "00000000",
   5364=> "01000000"
        & "00100000",
   5365=> "11111000"
        & "00100000",
   5366=> "00100000"
        & "00100000",
   5367=> "11111000"
        & "00000000",
   5368=> "01010000"
        & "00000000",
   5369=> "11111000"
        & "00100000",
   5370=> "00100000"
        & "00100000",
   5371=> "11111000"
        & "00000000",
   5372=> "00100000"
        & "01010000",
   5373=> "11111000"
        & "00100000",
   5374=> "00100000"
        & "00100000",
   5375=> "11111000"
        & "00000000",
   5376=> "00010000"
        & "00100000",
   5377=> "01110000"
        & "10001000",
   5378=> "10001000"
        & "10001000",
   5379=> "01110000"
        & "00000000",
   5380=> "01000000"
        & "00100000",
   5381=> "01110000"
        & "10001000",
   5382=> "10001000"
        & "10001000",
   5383=> "01110000"
        & "00000000",
   5384=> "01010000"
        & "00000000",
   5385=> "01110000"
        & "10001000",
   5386=> "10001000"
        & "10001000",
   5387=> "01110000"
        & "00000000",
   5388=> "00100000"
        & "01010000",
   5389=> "01110000"
        & "10001000",
   5390=> "10001000"
        & "10001000",
   5391=> "01110000"
        & "00000000",
   5392=> "00010000"
        & "00100000",
   5393=> "10001000"
        & "10001000",
   5394=> "10001000"
        & "10001000",
   5395=> "01110000"
        & "00000000",
   5396=> "01000000"
        & "00100000",
   5397=> "10001000"
        & "10001000",
   5398=> "10001000"
        & "10001000",
   5399=> "01110000"
        & "00000000",
   5400=> "01010000"
        & "00000000",
   5401=> "10001000"
        & "10001000",
   5402=> "10001000"
        & "10001000",
   5403=> "01110000"
        & "00000000",
   5404=> "00100000"
        & "01010000",
   5405=> "00000000"
        & "10001000",
   5406=> "10001000"
        & "10001000",
   5407=> "01110000"
        & "00000000",
   5408=> "00010000"
        & "00100000",
   5409=> "01110000"
        & "00001000",
   5410=> "01111000"
        & "10001000",
   5411=> "01111000"
        & "00000000",
   5412=> "01000000"
        & "00100000",
   5413=> "01110000"
        & "00001000",
   5414=> "01111000"
        & "10001000",
   5415=> "01111000"
        & "00000000",
   5416=> "01010000"
        & "00000000",
   5417=> "01110000"
        & "00001000",
   5418=> "01111000"
        & "10001000",
   5419=> "01111000"
        & "00000000",
   5420=> "00100000"
        & "01010000",
   5421=> "01110000"
        & "00001000",
   5422=> "01111000"
        & "10001000",
   5423=> "01111000"
        & "00000000",
   5424=> "00010000"
        & "00100000",
   5425=> "01111000"
        & "10000100",
   5426=> "11111100"
        & "10000000",
   5427=> "01111100"
        & "00000000",
   5428=> "00100000"
        & "00010000",
   5429=> "01111000"
        & "10000100",
   5430=> "11111100"
        & "10000000",
   5431=> "01111100"
        & "00000000",
   5432=> "01010000"
        & "00000000",
   5433=> "01111000"
        & "10000100",
   5434=> "11111100"
        & "10000000",
   5435=> "01111100"
        & "00000000",
   5436=> "00100000"
        & "01010000",
   5437=> "01111000"
        & "10000100",
   5438=> "11111100"
        & "10000000",
   5439=> "01111100"
        & "00000000",
   5440=> "00010000"
        & "00100000",
   5441=> "00000000"
        & "01100000",
   5442=> "00100000"
        & "00100000",
   5443=> "01110000"
        & "00000000",
   5444=> "01000000"
        & "00100000",
   5445=> "00000000"
        & "01100000",
   5446=> "00100000"
        & "00100000",
   5447=> "01110000"
        & "00000000",
   5448=> "00000000"
        & "01010000",
   5449=> "00000000"
        & "01100000",
   5450=> "00100000"
        & "00100000",
   5451=> "01110000"
        & "00000000",
   5452=> "00100000"
        & "01010000",
   5453=> "00000000"
        & "01100000",
   5454=> "00100000"
        & "00100000",
   5455=> "01110000"
        & "00000000",
   5456=> "00010000"
        & "00100000",
   5457=> "00000000"
        & "01110000",
   5458=> "10001000"
        & "10001000",
   5459=> "01110000"
        & "00000000",
   5460=> "01000000"
        & "00100000",
   5461=> "00000000"
        & "01110000",
   5462=> "10001000"
        & "10001000",
   5463=> "01110000"
        & "00000000",
   5464=> "00000000"
        & "01010000",
   5465=> "00000000"
        & "01110000",
   5466=> "10001000"
        & "10001000",
   5467=> "01110000"
        & "00000000",
   5468=> "00100000"
        & "01010000",
   5469=> "00000000"
        & "01110000",
   5470=> "10001000"
        & "10001000",
   5471=> "01110000"
        & "00000000",
   5472=> "00010000"
        & "00100000",
   5473=> "00000000"
        & "10001000",
   5474=> "10001000"
        & "10011000",
   5475=> "01101000"
        & "00000000",
   5476=> "01000000"
        & "00100000",
   5477=> "00000000"
        & "10001000",
   5478=> "10001000"
        & "10011000",
   5479=> "01101000"
        & "00000000",
   5480=> "00000000"
        & "01010000",
   5481=> "00000000"
        & "10001000",
   5482=> "10001000"
        & "10011000",
   5483=> "01101000"
        & "00000000",
   5484=> "00100000"
        & "01010000",
   5485=> "00000000"
        & "10001000",
   5486=> "10001000"
        & "10011000",
   5487=> "01101000"
        & "00000000",
   5488=> "01010000"
        & "00000000",
   5489=> "10001000"
        & "01010000",
   5490=> "00100000"
        & "00100000",
   5491=> "00100000"
        & "00000000",
   5492=> "01010000"
        & "00000000",
   5493=> "10001000"
        & "01010000",
   5494=> "00100000"
        & "01000000",
   5495=> "10000000"
        & "00000000",
   5496=> "00100000"
        & "00000000",
   5497=> "00100000"
        & "01000000",
   5498=> "10000000"
        & "10001000",
   5499=> "01110000"
        & "00000000",
   5500=> "00100000"
        & "00100000",
   5501=> "00000000"
        & "00100000",
   5502=> "00100000"
        & "00100000",
   5503=> "00100000"
        & "00000000",
   5504=> "00000000"
        & "00000000",
   5505=> "01001000"
        & "10010000",
   5506=> "01001000"
        & "00000000",
   5507=> "00000000"
        & "00000000",
   5508=> "00000000"
        & "00000000",
   5509=> "10010000"
        & "01001000",
   5510=> "10010000"
        & "00000000",
   5511=> "00000000"
        & "00000000",
   5512=> "10001000"
        & "00100010",
   5513=> "10001000"
        & "00100010",
   5514=> "10001000"
        & "00100010",
   5515=> "10001000"
        & "00100010",
   5516=> "10101010"
        & "01010101",
   5517=> "10101010"
        & "01010101",
   5518=> "10101010"
        & "01010101",
   5519=> "10101010"
        & "01010100",
   5520=> "11001100"
        & "11111111",
   5521=> "00110011"
        & "11001100",
   5522=> "11111111"
        & "00110011",
   5523=> "11001100"
        & "11111111",
   5524=> "00110000"
        & "00110000",
   5525=> "00110000"
        & "00110000",
   5526=> "00110000"
        & "00110000",
   5527=> "00110000"
        & "00110000",
   5528=> "00000000"
        & "00000000",
   5529=> "00000000"
        & "11111100",
   5530=> "11111100"
        & "00000000",
   5531=> "00000000"
        & "00000000",
   5532=> "00110000"
        & "00110000",
   5533=> "00110000"
        & "00111100",
   5534=> "00111100"
        & "00000000",
   5535=> "00000000"
        & "00000000",
   5536=> "00110000"
        & "00110000",
   5537=> "00110000"
        & "11110000",
   5538=> "11110000"
        & "00000000",
   5539=> "00000000"
        & "00000000",
   5540=> "00000000"
        & "00000000",
   5541=> "00000000"
        & "00111100",
   5542=> "00111100"
        & "00110000",
   5543=> "00110000"
        & "00110000",
   5544=> "00000000"
        & "00000000",
   5545=> "00000000"
        & "11110000",
   5546=> "11110000"
        & "00110000",
   5547=> "00110000"
        & "00110000",
   5548=> "00110000"
        & "00110000",
   5549=> "00110000"
        & "11110000",
   5550=> "11110000"
        & "00110000",
   5551=> "00110000"
        & "00110000",
   5552=> "00110000"
        & "00110000",
   5553=> "00110000"
        & "11111100",
   5554=> "11111100"
        & "00000000",
   5555=> "00000000"
        & "00000000",
   5556=> "00110000"
        & "00110000",
   5557=> "00110000"
        & "00111100",
   5558=> "00111100"
        & "00110000",
   5559=> "00110000"
        & "00110000",
   5560=> "00000000"
        & "00000000",
   5561=> "00000000"
        & "11111100",
   5562=> "11111100"
        & "00110000",
   5563=> "00110000"
        & "00110000",
   5564=> "00110000"
        & "00110000",
   5565=> "00110000"
        & "11111100",
   5566=> "11111100"
        & "00110000",
   5567=> "00110000"
        & "00110000",
   5568=> "00110000"
        & "00110000",
   5569=> "00110000"
        & "00110000",
   5570=> "00110000"
        & "00000000",
   5571=> "00000000"
        & "00000000",
   5572=> "00000000"
        & "00000000",
   5573=> "00000000"
        & "11110000",
   5574=> "11110000"
        & "00000000",
   5575=> "00000000"
        & "00000000",
   5576=> "00000000"
        & "00000000",
   5577=> "00000000"
        & "00111100",
   5578=> "00111100"
        & "00000000",
   5579=> "00000000"
        & "00000000",
   5580=> "00000000"
        & "00000000",
   5581=> "00000000"
        & "00110000",
   5582=> "00110000"
        & "00110000",
   5583=> "00110000"
        & "00110000",
   5584=> "11111100"
        & "10000100",
   5585=> "10000100"
        & "10000100",
   5586=> "10000100"
        & "10000100",
   5587=> "10000100"
        & "11111100",
   5588=> "11111100"
        & "11111100",
   5589=> "11001100"
        & "11001100",
   5590=> "11001100"
        & "11001100",
   5591=> "11111100"
        & "11111100",
   5592=> "11111100"
        & "11111100",
   5593=> "11111100"
        & "11111100",
   5594=> "11111100"
        & "11111100",
   5595=> "11111100"
        & "11111100",
   5596=> "11111100"
        & "11111100",
   5597=> "11111100"
        & "11111100",
   5598=> "00000000"
        & "00000000",
   5599=> "00000000"
        & "00000000",
   5600=> "11100000"
        & "11100000",
   5601=> "11100000"
        & "11100000",
   5602=> "11100000"
        & "11100000",
   5603=> "11100000"
        & "11100000",
   5604=> "00011100"
        & "00011100",
   5605=> "00011100"
        & "00011100",
   5606=> "00011100"
        & "00011100",
   5607=> "00011100"
        & "00011100",
   5608=> "00000000"
        & "00000000",
   5609=> "00000000"
        & "00000000",
   5610=> "11111100"
        & "11111100",
   5611=> "11111100"
        & "11111100",
   5612=> "00000000"
        & "00000000",
   5613=> "01101000"
        & "10010000",
   5614=> "10010000"
        & "10010000",
   5615=> "01101000"
        & "00000000",
   5616=> "00110000"
        & "01001000",
   5617=> "01001000"
        & "01110000",
   5618=> "01001000"
        & "01101000",
   5619=> "01010000"
        & "00000000",
   5620=> "00000000"
        & "11111000",
   5621=> "10000000"
        & "10000000",
   5622=> "10000000"
        & "10000000",
   5623=> "10000000"
        & "00000000",
   5624=> "00000000"
        & "01000000",
   5625=> "10101000"
        & "00010000",
   5626=> "00010000"
        & "00010000",
   5627=> "00010000"
        & "00000000",
   5628=> "00100000"
        & "00100000",
   5629=> "01010000"
        & "01010000",
   5630=> "10001000"
        & "10001000",
   5631=> "11111000"
        & "00000000",
   5632=> "01110000"
        & "10001000",
   5633=> "01100000"
        & "00010000",
   5634=> "01110000"
        & "10001000",
   5635=> "01110000"
        & "00000000",
   5636=> "00000000"
        & "00000000",
   5637=> "01111000"
        & "10000000",
   5638=> "11111000"
        & "10000000",
   5639=> "01111000"
        & "00000000",
   5640=> "00100000"
        & "00011000",
   5641=> "00100000"
        & "01000000",
   5642=> "00110000"
        & "00001000",
   5643=> "01110000"
        & "00000000",
   5644=> "01110000"
        & "10001000",
   5645=> "10001000"
        & "11111000",
   5646=> "10001000"
        & "10001000",
   5647=> "01110000"
        & "00000000",
   5648=> "00000000"
        & "00000000",
   5649=> "11000000"
        & "01000000",
   5650=> "01000000"
        & "01010000",
   5651=> "00100000"
        & "00000000",
   5652=> "00100000"
        & "00100000",
   5653=> "01010000"
        & "01010000",
   5654=> "10001000"
        & "10001000",
   5655=> "10001000"
        & "00000000",
   5656=> "00000000"
        & "11000000",
   5657=> "00100000"
        & "00100000",
   5658=> "01010000"
        & "01001000",
   5659=> "10001000"
        & "00000000",
   5660=> "00000000"
        & "00000000",
   5661=> "10010000"
        & "10000000",
   5662=> "10010000"
        & "11111000",
   5663=> "10000000"
        & "00000000",
   5664=> "00000000"
        & "11111000",
   5665=> "10001000"
        & "10001000",
   5666=> "10001000"
        & "10001000",
   5667=> "10001000"
        & "00000000",
   5668=> "00000000"
        & "00000000",
   5669=> "00000000"
        & "11111000",
   5670=> "01010000"
        & "01010000",
   5671=> "01010000"
        & "00000000",
   5672=> "11111100"
        & "01000000",
   5673=> "00100000"
        & "00010000",
   5674=> "00100000"
        & "01000000",
   5675=> "11111000"
        & "00000000",
   5676=> "00000000"
        & "00000000",
   5677=> "01111000"
        & "10010000",
   5678=> "10010000"
        & "10010000",
   5679=> "01100000"
        & "00000000",
   5680=> "00000000"
        & "00000000",
   5681=> "01111000"
        & "10100000",
   5682=> "00100000"
        & "00100000",
   5683=> "00011000"
        & "00000000",
   5684=> "00100000"
        & "00100000",
   5685=> "01110000"
        & "10101000",
   5686=> "01110000"
        & "00100000",
   5687=> "00100000"
        & "00000000",
   5688=> "10000000"
        & "01001000",
   5689=> "01010000"
        & "00100000",
   5690=> "01010000"
        & "10010000",
   5691=> "00001000"
        & "00000000",
   5692=> "00000000"
        & "01110000",
   5693=> "10001000"
        & "10001000",
   5694=> "10001000"
        & "01010000",
   5695=> "11011000"
        & "00000000",
   5696=> "00000000"
        & "11111000",
   5697=> "00000000"
        & "11111000",
   5698=> "00000000"
        & "11111000",
   5699=> "00000000"
        & "00000000",
   5700=> "00000000"
        & "00100000",
   5701=> "00100000"
        & "11111000",
   5702=> "00100000"
        & "00100000",
   5703=> "11111000"
        & "00000000",
   5704=> "11000000"
        & "00110000",
   5705=> "00001000"
        & "00110000",
   5706=> "11000000"
        & "00000000",
   5707=> "11111000"
        & "00000000",
   5708=> "00011000"
        & "01100000",
   5709=> "10000000"
        & "01100000",
   5710=> "00011000"
        & "00000000",
   5711=> "11111000"
        & "00000000",
   5712=> "00000000"
        & "00100000",
   5713=> "00000000"
        & "11111000",
   5714=> "00000000"
        & "00100000",
   5715=> "00000000"
        & "00000000",
   5716=> "00110000"
        & "01001000",
   5717=> "00110000"
        & "00000000",
   5718=> "00000000"
        & "00000000",
   5719=> "00000000"
        & "00000000",
   5720=> "00000000"
        & "00011000",
   5721=> "00010000"
        & "00010000",
   5722=> "10010000"
        & "01010000",
   5723=> "00100000"
        & "00000000",
   5724=> "01100000"
        & "00010000",
   5725=> "00100000"
        & "01110000",
   5726=> "00000000"
        & "00000000",
   5727=> "00000000"
        & "00000000",
   5728=> "01110000"
        & "10001000",
   5729=> "10001000"
        & "10010000",
   5730=> "10001000"
        & "10001000",
   5731=> "10001000"
        & "10110000",
   5732=> "00000000"
        & "00100000",
   5733=> "01110000"
        & "10100000",
   5734=> "10100000"
        & "01110000",
   5735=> "00100000"
        & "00000000",
   5736=> "00111100"
        & "01010000",
   5737=> "10010000"
        & "11111100",
   5738=> "10010000"
        & "10010000",
   5739=> "10011100"
        & "00000000",
   5740=> "01111100"
        & "10010000",
   5741=> "10010000"
        & "10011100",
   5742=> "10010000"
        & "10010000",
   5743=> "01111100"
        & "00000000",
   5744=> "01110000"
        & "10001000",
   5745=> "10000000"
        & "11110000",
   5746=> "01000000"
        & "01000000",
   5747=> "11111000"
        & "00000000",
   5748=> "10001000"
        & "10001000",
   5749=> "01010000"
        & "11111000",
   5750=> "00100000"
        & "11111000",
   5751=> "00100000"
        & "00000000",
   5752=> "00010000"
        & "00101000",
   5753=> "00100000"
        & "00100000",
   5754=> "00100000"
        & "10100000",
   5755=> "01000000"
        & "00000000",
   5756=> "11111000"
        & "10000000",
   5757=> "10000000"
        & "11110000",
   5758=> "10001000"
        & "10001000",
   5759=> "11110000"
        & "00000000",
   5760=> "11110000"
        & "01010000",
   5761=> "01010000"
        & "10010000",
   5762=> "10010000"
        & "11111000",
   5763=> "10001000"
        & "00000000",
   5764=> "10101000"
        & "10101000",
   5765=> "01110000"
        & "10101000",
   5766=> "10101000"
        & "10101000",
   5767=> "10101000"
        & "00000000",
   5768=> "01110000"
        & "10001000",
   5769=> "00001000"
        & "00110000",
   5770=> "00001000"
        & "10001000",
   5771=> "01110000"
        & "00000000",
   5772=> "10001000"
        & "10001000",
   5773=> "11001000"
        & "10101000",
   5774=> "10011000"
        & "10001000",
   5775=> "10001000"
        & "00000000",
   5776=> "01010000"
        & "00100000",
   5777=> "10001000"
        & "11001000",
   5778=> "10101000"
        & "10011000",
   5779=> "10001000"
        & "00000000",
   5780=> "01111000"
        & "01001000",
   5781=> "01001000"
        & "01001000",
   5782=> "01001000"
        & "01001000",
   5783=> "11001000"
        & "00000000",
   5784=> "10001000"
        & "10001000",
   5785=> "10001000"
        & "10001000",
   5786=> "10001000"
        & "11111000",
   5787=> "00001000"
        & "00000000",
   5788=> "10001000"
        & "10001000",
   5789=> "10001000"
        & "01111000",
   5790=> "00001000"
        & "00001000",
   5791=> "00001000"
        & "00000000",
   5792=> "10101000"
        & "10101000",
   5793=> "10101000"
        & "10101000",
   5794=> "10101000"
        & "10101000",
   5795=> "11111000"
        & "00000000",
   5796=> "10101000"
        & "10101000",
   5797=> "10101000"
        & "10101000",
   5798=> "10101000"
        & "11111000",
   5799=> "00001000"
        & "00000000",
   5800=> "11000000"
        & "01000000",
   5801=> "01000000"
        & "01110000",
   5802=> "01001000"
        & "01001000",
   5803=> "01110000"
        & "00000000",
   5804=> "10001000"
        & "10001000",
   5805=> "10001000"
        & "11101000",
   5806=> "10011000"
        & "10011000",
   5807=> "11101000"
        & "00000000",
   5808=> "10000000"
        & "10000000",
   5809=> "10000000"
        & "11110000",
   5810=> "10001000"
        & "10001000",
   5811=> "11110000"
        & "00000000",
   5812=> "01110000"
        & "10001000",
   5813=> "00001000"
        & "01111000",
   5814=> "00001000"
        & "10001000",
   5815=> "01110000"
        & "00000000",
   5816=> "10010000"
        & "10101000",
   5817=> "10101000"
        & "11101000",
   5818=> "10101000"
        & "10101000",
   5819=> "10010000"
        & "00000000",
   5820=> "01111000"
        & "10001000",
   5821=> "10001000"
        & "01111000",
   5822=> "01001000"
        & "10001000",
   5823=> "10001000"
        & "00000000",
   
   -- Hello World\0
   5824=> x"48"
        & x"65",
   5825=> x"6C"
        & x"6C",
   5826=> x"6F"
        & x"20",
   5827=> x"57"
        & x"6F",
   5828=> x"72"
        & x"6C",
   5829=> x"64"
        & x"00",

 
 others => x"0000"
 );
begin
   process(CLK)
	begin 
		if (CLK'event AND CLK='1') then
			DOUT2 <= memoire(to_integer(unsigned(AD2)));
		end if;
	end process;

	process(CLK)
	begin 
		if (CLK'event AND CLK='1') then
			if ((CE1='1') AND (OE1='1')) then 
				DOUT1<=memoire(to_integer(unsigned(AD1)));
			else 
				DOUT1<=(others =>'0');
			end if;		
		end if;
	end process;
	
	process (CLK)
	begin
	  IF (CLK'event AND CLK='1') then
			if ((CE1='1') AND (WE1='1')) then 
				memoire(to_integer(unsigned(AD1)))<=DIN1;
			end if;
		  end if;
	end process;
	
end Behavioral;

