----------------------------------------------------------------------------------
--
-- File retrieved, on 07/02/2010, from :
-- http://sebastien-viardot.imag.fr/Enseignements/Archi1A2s/sources/ROMPROG.vhd
--
-- Slightly altered to get rid of vendor-specific packages and adjust formatting
-- Now auto-filled by asrom script
--
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROMPROG is
  Port ( AD : in  STD_LOGIC_VECTOR (12 downto 0);
         D : out  STD_LOGIC_VECTOR (15 downto 0);
         CLK : in STD_LOGIC);
end ROMPROG;

architecture Behavioral of ROMPROG is
  constant low_address: natural := 0;
  constant high_address: natural := 8192;
  subtype octet is std_logic_vector( 15 downto 0 );
  type zone_memoire is
    array (natural range low_address to high_address-1) of octet;
  constant m: zone_memoire:= (
    0=>x"FFF7",	-- 1111111111110111  liw	r7, IRQ_mask
    1=>x"2000",	-- 0010000000000000  
    2=>x"F8C0",	-- 1111100011000000  bai	-, os_init
    3=>x"0100",	-- 0000000100000000  
   16=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_ack
   17=>x"2002",	-- 0010000000000010  
   18=>x"D001",	-- 1101000000000001  lw	r1, r0
   19=>x"F54A",	-- 1111010101001010  bspl	r2, r1, 5
   20=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_error
   21=>x"0050",	-- 0000000001010000  
   22=>x"F4CA",	-- 1111010011001010  bspl	r2, r1, 3
   23=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_kbd
   24=>x"0060",	-- 0000000001100000  
   25=>x"F40A",	-- 1111010000001010  bspl	r2, r1, 0
   26=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_tmr
   27=>x"0040",	-- 0000000001000000  
   28=>x"D201",	-- 1101001000000001  sw	r1, r0
   29=>x"FFFE",	-- 1111111111111110  reti
   64=>x"263F",	-- 0010011000111111  not r7, r7
   65=>x"D7C0",	-- 1101011111000000  out	r7
   66=>x"E383",	-- 1110001110000011  ba	-, r6
   80=>x"25FF",	-- 0010010111111111  xor	r7, r7, r7
   81=>x"D7C0",	-- 1101011111000000  out	r7
   82=>x"E383",	-- 1110001110000011  ba	-, r6
   96=>x"FFF2",	-- 1111111111110010  liw	r2, PS2_rx
   97=>x"2004",	-- 0010000000000100  
   98=>x"D012",	-- 1101000000010010  lw	r2, r2
   99=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map + 8
  100=>x"1808",	-- 0001100000001000  
  101=>x"D01B",	-- 1101000000011011  lw	r3, r3
  102=>x"1EBF",	-- 0001111010111111  mixll	r7, r7, r2
  103=>x"C784",	-- 1100011110000100  li	r4, 0xF0
  104=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  105=>x"8B20",	-- 1000101100100000  brieq	r4, int_kbd.release
  106=>x"C704",	-- 1100011100000100  li	r4, 0xE0
  107=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  108=>x"88E0",	-- 1000100011100000  brieq	r4, int_kbd.extended
  109=>x"FFF5",	-- 1111111111110101  liw	r5, paper_keys - 1
  110=>x"16BF",	-- 0001011010111111  
  111=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  112=>x"80E0",	-- 1000000011100000  brieq	r4, $+3
  113=>x"FFF5",	-- 1111111111110101  liw	r5, paper_keys + 11 - 1
  114=>x"16CA",	-- 0001011011001010  
  115=>x"042D",	-- 0000010000101101  inc	r5, r5
  116=>x"D02C",	-- 1101000000101100  lw	r4, r5
  117=>x"8560",	-- 1000010101100000  brieq	r4, scan_code_mismatch
  118=>x"6E24",	-- 0110111000100100  shr	r4, r4, 7
  119=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  120=>x"BEE4",	-- 1011111011100100  brine	r4, scan_code_loop
  121=>x"D02A",	-- 1101000000101010  lw	r2, r5
  122=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  123=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  124=>x"741B",	-- 0111010000011011  shr	r3, r3, 10
  125=>x"C00D",	-- 1100000000001101  li	r5, 1
  126=>x"0612",	-- 0000011000010010  dec	r2, r2
  127=>x"3AAA",	-- 0011101010101010  rrl	r2, r5, r2
  128=>x"FFF5",	-- 1111111111110101  liw	r5, key_press_map
  129=>x"1800",	-- 0001100000000000  
  130=>x"08ED",	-- 0000100011101101  add	r5, r5, r3
  131=>x"D02B",	-- 1101000000101011  lw	r3, r5
  132=>x"80E4",	-- 1000000011100100  brine	r4, scan_code_release
  133=>x"229B",	-- 0010001010011011  or	r3, r3, r2
  134=>x"80C3",	-- 1000000011000011  bri	-, scan_code_notify
  135=>x"2612",	-- 0010011000010010  not	r2, r2
  136=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  137=>x"D22B",	-- 1101001000101011  sw	r3, r5
  138=>x"C003",	-- 1100000000000011  li	r3, 0
  139=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  140=>x"1808",	-- 0001100000001000  
  141=>x"D223",	-- 1101001000100011  sw	r3, r4
  142=>x"E383",	-- 1110001110000011  ba	-, r6
  143=>x"C014",	-- 1100000000010100  li	r4, 2
  144=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  145=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  146=>x"1808",	-- 0001100000001000  
  147=>x"D223",	-- 1101001000100011  sw	r3, r4
  148=>x"E383",	-- 1110001110000011  ba	-, r6
  149=>x"C00C",	-- 1100000000001100  li	r4, 1
  150=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  151=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  152=>x"1808",	-- 0001100000001000  
  153=>x"D223",	-- 1101001000100011  sw	r3, r4
  154=>x"E383",	-- 1110001110000011  ba	-, r6
  256=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_mask
  257=>x"2000",	-- 0010000000000000  
  258=>x"C0C9",	-- 1100000011001001  li	r1, 0x19
  259=>x"D201",	-- 1101001000000001  sw	r1, r0
  260=>x"0400",	-- 0000010000000000  inc	r0, r0
  261=>x"CFF9",	-- 1100111111111001  li	r1, -1
  262=>x"D201",	-- 1101001000000001  sw	r1, r0
  263=>x"C03A",	-- 1100000000111010  li	r2, 7
  264=>x"0880",	-- 0000100010000000  add	r0, r0, r2
  265=>x"C0EA",	-- 1100000011101010  li	r2, 0x1D
  266=>x"D202",	-- 1101001000000010  sw	r2, r0
  267=>x"0400",	-- 0000010000000000  inc	r0, r0
  268=>x"C07A",	-- 1100000001111010  li	r2, 15
  269=>x"D202",	-- 1101001000000010  sw	r2, r0
  270=>x"FFF0",	-- 1111111111110000  liw	r0, key_press_map
  271=>x"1800",	-- 0001100000000000  
  272=>x"C001",	-- 1100000000000001  li	r1, 0
  273=>x"C042",	-- 1100000001000010  li	r2, 8
  274=>x"D201",	-- 1101001000000001  sw	r1, r0
  275=>x"0400",	-- 0000010000000000  inc	r0, r0
  276=>x"0612",	-- 0000011000010010  dec	r2, r2
  277=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  278=>x"C0F3",	-- 1100000011110011  li	r3, 30
  279=>x"CFFA",	-- 1100111111111010  li	r2, -1
  280=>x"D21A",	-- 1101001000011010  sw	r2, r3
  281=>x"8083",	-- 1000000010000011  bri	-, PaperGameStart
  282=>x"8003",	-- 1000000000000011  bri	-, PaperMenuLoop
  283=>x"FFF0",	-- 1111111111110000  liw	r0, paper_dir
  284=>x"1732",	-- 0001011100110010  
  285=>x"C001",	-- 1100000000000001  li	r1, 0
  286=>x"D201",	-- 1101001000000001  sw	r1, r0
  287=>x"0400",	-- 0000010000000000  inc	r0, r0
  288=>x"C4C1",	-- 1100010011000001  li	r1, 152
  289=>x"D201",	-- 1101001000000001  sw	r1, r0
  290=>x"0400",	-- 0000010000000000  inc	r0, r0
  291=>x"C001",	-- 1100000000000001  li	r1, 0
  292=>x"D201",	-- 1101001000000001  sw	r1, r0
  293=>x"0400",	-- 0000010000000000  inc	r0, r0
  294=>x"C401",	-- 1100010000000001  li	r1, 128
  295=>x"D201",	-- 1101001000000001  sw	r1, r0
  296=>x"0400",	-- 0000010000000000  inc	r0, r0
  297=>x"C001",	-- 1100000000000001  li	r1, 0
  298=>x"D201",	-- 1101001000000001  sw	r1, r0
  299=>x"0400",	-- 0000010000000000  inc	r0, r0
  300=>x"C0A1",	-- 1100000010100001  li	r1, 20
  301=>x"D201",	-- 1101001000000001  sw	r1, r0
  302=>x"0400",	-- 0000010000000000  inc	r0, r0
  303=>x"C029",	-- 1100000000101001  li	r1, 5
  304=>x"D201",	-- 1101001000000001  sw	r1, r0
  305=>x"0400",	-- 0000010000000000  inc	r0, r0
  306=>x"C000",	-- 1100000000000000  li	r0, 0
  307=>x"CFF9",	-- 1100111111111001  li	r1, -1
  308=>x"C0A2",	-- 1100000010100010  li	r2, 20
  309=>x"D201",	-- 1101001000000001  sw	r1, r0
  310=>x"0400",	-- 0000010000000000  inc	r0, r0
  311=>x"0612",	-- 0000011000010010  dec	r2, r2
  312=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  313=>x"C001",	-- 1100000000000001  li	r1, 0
  314=>x"FFF2",	-- 1111111111110010  liw	r2, 18*20
  315=>x"0168",	-- 0000000101101000  
  316=>x"D201",	-- 1101001000000001  sw	r1, r0
  317=>x"0400",	-- 0000010000000000  inc	r0, r0
  318=>x"0612",	-- 0000011000010010  dec	r2, r2
  319=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  320=>x"CFF9",	-- 1100111111111001  li	r1, -1
  321=>x"C0A2",	-- 1100000010100010  li	r2, 20
  322=>x"D201",	-- 1101001000000001  sw	r1, r0
  323=>x"0400",	-- 0000010000000000  inc	r0, r0
  324=>x"0612",	-- 0000011000010010  dec	r2, r2
  325=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  326=>x"C020",	-- 1100000000100000  li	r0, 4
  327=>x"C029",	-- 1100000000101001  li	r1, 5
  328=>x"FFF2",	-- 1111111111110010  liw	r2, paper_title
  329=>x"173A",	-- 0001011100111010  
  330=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  331=>x"0215",	-- 0000001000010101  
  332=>x"C788",	-- 1100011110001000  li	r0, 241
  333=>x"C009",	-- 1100000000001001  li	r1, 1
  334=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud
  335=>x"1720",	-- 0001011100100000  
  336=>x"C043",	-- 1100000001000011  li	r3, 8
  337=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  338=>x"02BF",	-- 0000001010111111  
  339=>x"C0F8",	-- 1100000011111000  li	r0, 31
  340=>x"C009",	-- 1100000000001001  li	r1, 1
  341=>x"C3DA",	-- 1100001111011010  li	r2, 123
  342=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum
  343=>x"0244",	-- 0000001001000100  
  344=>x"C120",	-- 1100000100100000  li	r0, 36
  345=>x"C009",	-- 1100000000001001  li	r1, 1
  346=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  347=>x"1741",	-- 0001011101000001  
  348=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  349=>x"0215",	-- 0000001000010101  
  350=>x"C788",	-- 1100011110001000  li	r0, 241
  351=>x"C051",	-- 1100000001010001  li	r1, 10
  352=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud + 4
  353=>x"1724",	-- 0001011100100100  
  354=>x"C043",	-- 1100000001000011  li	r3, 8
  355=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  356=>x"02BF",	-- 0000001010111111  
  357=>x"C0F8",	-- 1100000011111000  li	r0, 31
  358=>x"C051",	-- 1100000001010001  li	r1, 10
  359=>x"C16A",	-- 1100000101101010  li	r2, 45
  360=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum
  361=>x"0244",	-- 0000001001000100  
  362=>x"C120",	-- 1100000100100000  li	r0, 36
  363=>x"C051",	-- 1100000001010001  li	r1, 10
  364=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  365=>x"1741",	-- 0001011101000001  
  366=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  367=>x"0215",	-- 0000001000010101  
  368=>x"FFF0",	-- 1111111111110000  liw	r0, 20*20
  369=>x"0190",	-- 0000000110010000  
  370=>x"C001",	-- 1100000000000001  li	r1, 0
  371=>x"FFF2",	-- 1111111111110010  liw	r2, 220*20
  372=>x"1130",	-- 0001000100110000  
  373=>x"D201",	-- 1101001000000001  sw	r1, r0
  374=>x"0400",	-- 0000010000000000  inc	r0, r0
  375=>x"0612",	-- 0000011000010010  dec	r2, r2
  376=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  377=>x"FFF5",	-- 1111111111110101  liw	r5, paper_tilemap
  378=>x"1780",	-- 0001011110000000  
  379=>x"D02C",	-- 1101000000101100  lw	r4, r5
  380=>x"042D",	-- 0000010000101101  inc	r5, r5
  381=>x"8620",	-- 1000011000100000  brieq	r4, PaperGameTileSkip
  382=>x"063F",	-- 0000011000111111  dec	r7, r7
  383=>x"D23D",	-- 1101001000111101  sw	r5, r7
  384=>x"FFF3",	-- 1111111111110011  liw	r3, paper_tilemap
  385=>x"1780",	-- 0001011110000000  
  386=>x"0AEB",	-- 0000101011101011  sub	r3, r5, r3
  387=>x"6E20",	-- 0110111000100000  shr	r0, r4, 7
  388=>x"6219",	-- 0110001000011001  shr	r1, r3, 1
  389=>x"4609",	-- 0100011000001001  shl	r1, r1, 3
  390=>x"C00B",	-- 1100000000001011  li	r3, 1
  391=>x"FB06",	-- 1111101100000110  bailne	r0, r6, put_tile
  392=>x"01CD",	-- 0000000111001101  
  393=>x"4E24",	-- 0100111000100100  shl	r4, r4, 7
  394=>x"6E24",	-- 0110111000100100  shr	r4, r4, 7
  395=>x"C013",	-- 1100000000010011  li	r3, 2
  396=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_tile
  397=>x"01CD",	-- 0000000111001101  
  398=>x"0624",	-- 0000011000100100  dec	r4, r4
  399=>x"BF24",	-- 1011111100100100  brine	r4, PaperGameSegmentLoop
  400=>x"C003",	-- 1100000000000011  li	r3, 0
  401=>x"FB06",	-- 1111101100000110  bailne	r0, r6, put_tile
  402=>x"01CD",	-- 0000000111001101  
  403=>x"D03D",	-- 1101000000111101  lw	r5, r7
  404=>x"043F",	-- 0000010000111111  inc	r7, r7
  405=>x"FFF4",	-- 1111111111110100  liw r4, paper_tilemap + 125
  406=>x"17FD",	-- 0001011111111101  
  407=>x"0B2C",	-- 0000101100101100  sub	r4, r5, r4
  408=>x"B8E5",	-- 1011100011100101  brilt	r4, PaperGameTileLoop
  409=>x"FFF3",	-- 1111111111110011  liw	r3, paper_dir
  410=>x"1732",	-- 0001011100110010  
  411=>x"D01C",	-- 1101000000011100  lw	r4, r3
  412=>x"041B",	-- 0000010000011011  inc	r3, r3
  413=>x"D018",	-- 1101000000011000  lw	r0, r3
  414=>x"FFF2",	-- 1111111111110010  liw	r2, paper_sprites
  415=>x"16D0",	-- 0001011011010000  
  416=>x"4624",	-- 0100011000100100  shl	r4, r4, 3
  417=>x"0912",	-- 0000100100010010  add	r2, r2, r4
  418=>x"C161",	-- 1100000101100001  li	r1, 44
  419=>x"C083",	-- 1100000010000011  li	r3, 16
  420=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_16
  421=>x"0273",	-- 0000001001110011  
  422=>x"C02A",	-- 1100000000101010  li	r2, 5
  423=>x"C003",	-- 1100000000000011  li	r3, 0
  424=>x"061B",	-- 0000011000011011  dec	r3, r3
  425=>x"BFDC",	-- 1011111111011100  brine	r3, $-1
  426=>x"0612",	-- 0000011000010010  dec	r2, r2
  427=>x"BF14",	-- 1011111100010100  brine	r2, $-4
  428=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  429=>x"1800",	-- 0001100000000000  
  430=>x"D01B",	-- 1101000000011011  lw	r3, r3
  431=>x"BF58",	-- 1011111101011000  brieq	r3, PaperGameLoop
  432=>x"F7DC",	-- 1111011111011100  bspl	r4, r3, 15
  433=>x"86E4",	-- 1000011011100100  brine	r4, PaperGameQuit
  434=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  435=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveUp
  436=>x"F49C",	-- 1111010010011100  bspl	r4, r3, 2
  437=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveDOWN
  438=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  439=>x"82A0",	-- 1000001010100000  brieq	r4, PaperNoMoveLEFT
  440=>x"FFF2",	-- 1111111111110010  liw	r2, paper_dir
  441=>x"1732",	-- 0001011100110010  
  442=>x"C010",	-- 1100000000010000  li	r0, 2
  443=>x"D210",	-- 1101001000010000  sw	r0, r2
  444=>x"0412",	-- 0000010000010010  inc	r2, r2
  445=>x"D010",	-- 1101000000010000  lw	r0, r2
  446=>x"80C0",	-- 1000000011000000  brieq	r0, $+3
  447=>x"0600",	-- 0000011000000000  dec	r0, r0
  448=>x"D210",	-- 1101001000010000  sw	r0, r2
  449=>x"F4DC",	-- 1111010011011100  bspl	r4, r3, 3
  450=>x"8260",	-- 1000001001100000  brieq	r4, PaperNoMoveRIGHT
  451=>x"FFF2",	-- 1111111111110010  liw	r2, paper_dir
  452=>x"1732",	-- 0001011100110010  
  453=>x"C008",	-- 1100000000001000  li	r0, 1
  454=>x"D210",	-- 1101001000010000  sw	r0, r2
  455=>x"0412",	-- 0000010000010010  inc	r2, r2
  456=>x"D010",	-- 1101000000010000  lw	r0, r2
  457=>x"0400",	-- 0000010000000000  inc	r0, r0
  458=>x"D210",	-- 1101001000010000  sw	r0, r2
  459=>x"A943",	-- 1010100101000011  bri	-, PaperGameRedrawContent
  460=>x"FFFF",	-- 1111111111111111  reset
  461=>x"063F",	-- 0000011000111111  dec	r7, r7
  462=>x"D23E",	-- 1101001000111110  sw	r6, r7
  463=>x"063F",	-- 0000011000111111  dec	r7, r7
  464=>x"D238",	-- 1101001000111000  sw	r0, r7
  465=>x"063F",	-- 0000011000111111  dec	r7, r7
  466=>x"D239",	-- 1101001000111001  sw	r1, r7
  467=>x"063F",	-- 0000011000111111  dec	r7, r7
  468=>x"D23C",	-- 1101001000111100  sw	r4, r7
  469=>x"FFF2",	-- 1111111111110010  liw	r2, paper_tiles
  470=>x"1730",	-- 0001011100110000  
  471=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  472=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  473=>x"C043",	-- 1100000001000011  li	r3, 8
  474=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  475=>x"0299",	-- 0000001010011001  
  476=>x"D03C",	-- 1101000000111100  lw	r4, r7
  477=>x"043F",	-- 0000010000111111  inc	r7, r7
  478=>x"D039",	-- 1101000000111001  lw	r1, r7
  479=>x"043F",	-- 0000010000111111  inc	r7, r7
  480=>x"D038",	-- 1101000000111000  lw	r0, r7
  481=>x"043F",	-- 0000010000111111  inc	r7, r7
  482=>x"0400",	-- 0000010000000000  inc	r0, r0
  483=>x"D03E",	-- 1101000000111110  lw	r6, r7
  484=>x"043F",	-- 0000010000111111  inc	r7, r7
  485=>x"E383",	-- 1110001110000011  ba	-, r6
  486=>x"C750",	-- 1100011101010000  li	r0, 234
  487=>x"C1C2",	-- 1100000111000010  li	r2, 56
  488=>x"FAC6",	-- 1111101011000110  bail	-, r6, div_16_16
  489=>x"01FE",	-- 0000000111111110  
  490=>x"C448",	-- 1100010001001000  li	r0, 137
  491=>x"C472",	-- 1100010001110010  li	r2, 142
  492=>x"FAC6",	-- 1111101011000110  bail	-, r6, mult_16_16
  493=>x"01F2",	-- 0000000111110010  
  494=>x"C03A",	-- 1100000000111010  li r2, 7
  495=>x"FAC6",	-- 1111101011000110  bail	-, r6, fact_16
  496=>x"0209",	-- 0000001000001001  
  497=>x"FFFF",	-- 1111111111111111  reset
  498=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  499=>x"2524",	-- 0010010100100100  xor	r4, r4, r4
  500=>x"C085",	-- 1100000010000101  li	r5, 16
  501=>x"0849",	-- 0000100001001001  add	r1, r1, r1
  502=>x"0C00",	-- 0000110000000000  adc	r0, r0, r0
  503=>x"0EDB",	-- 0000111011011011  sbc	r3, r3, r3
  504=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  505=>x"08C9",	-- 0000100011001001  add	r1, r1, r3
  506=>x"0D00",	-- 0000110100000000  adc	r0, r0, r4
  507=>x"062D",	-- 0000011000101101  dec	r5, r5
  508=>x"BE6C",	-- 1011111001101100  brine	r5, mult_16_16.loop
  509=>x"E383",	-- 1110001110000011  ba	-, r6
  510=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  511=>x"C084",	-- 1100000010000100  li	r4, 16
  512=>x"0800",	-- 0000100000000000  add	r0, r0, r0
  513=>x"0C49",	-- 0000110001001001  adc	r1, r1, r1
  514=>x"0A8B",	-- 0000101010001011  sub	r3, r1, r2
  515=>x"80DD",	-- 1000000011011101  brilt	r3, div_16_16.skip
  516=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  517=>x"0400",	-- 0000010000000000  inc	r0, r0
  518=>x"0624",	-- 0000011000100100  dec	r4, r4
  519=>x"BE64",	-- 1011111001100100  brine	r4, div_16_16.loop
  520=>x"E383",	-- 1110001110000011  ba	-, r6
  521=>x"2400",	-- 0010010000000000  xor	r0, r0, r0
  522=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  523=>x"8250",	-- 1000001001010000  brieq	r2, fact_16.end
  524=>x"0409",	-- 0000010000001001  inc	r1, r1
  525=>x"1008",	-- 0001000000001000  mova	r0, r1
  526=>x"FAC6",	-- 1111101011000110  bail	-, r6, mult_16_16
  527=>x"01F2",	-- 0000000111110010  
  528=>x"8104",	-- 1000000100000100  brine	r0, fact_16.overflow
  529=>x"01F2",	-- 0000000111110010  
  530=>x"0612",	-- 0000011000010010  dec	r2, r2
  531=>x"BE94",	-- 1011111010010100  brine	r2, fact_16.loop
  532=>x"E383",	-- 1110001110000011  ba	-, r6
  533=>x"063F",	-- 0000011000111111  dec	r7, r7
  534=>x"D23E",	-- 1101001000111110  sw	r6, r7
  535=>x"D013",	-- 1101000000010011  lw	r3, r2
  536=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  537=>x"84D8",	-- 1000010011011000  brieq	r3, puts.end
  538=>x"063F",	-- 0000011000111111  dec	r7, r7
  539=>x"D23A",	-- 1101001000111010  sw	r2, r7
  540=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  541=>x"022F",	-- 0000001000101111  
  542=>x"D03A",	-- 1101000000111010  lw	r2, r7
  543=>x"043F",	-- 0000010000111111  inc	r7, r7
  544=>x"D013",	-- 1101000000010011  lw	r3, r2
  545=>x"4E1B",	-- 0100111000011011  shl	r3, r3, 7
  546=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  547=>x"8258",	-- 1000001001011000  brieq	r3, puts.end
  548=>x"063F",	-- 0000011000111111  dec	r7, r7
  549=>x"D23A",	-- 1101001000111010  sw	r2, r7
  550=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  551=>x"022F",	-- 0000001000101111  
  552=>x"D03A",	-- 1101000000111010  lw	r2, r7
  553=>x"043F",	-- 0000010000111111  inc	r7, r7
  554=>x"0412",	-- 0000010000010010  inc	r2, r2
  555=>x"BB03",	-- 1011101100000011  bri	-, puts.loop
  556=>x"D03E",	-- 1101000000111110  lw	r6, r7
  557=>x"043F",	-- 0000010000111111  inc	r7, r7
  558=>x"E383",	-- 1110001110000011  ba	-, r6
  559=>x"063F",	-- 0000011000111111  dec	r7, r7
  560=>x"D23E",	-- 1101001000111110  sw	r6, r7
  561=>x"063F",	-- 0000011000111111  dec	r7, r7
  562=>x"D238",	-- 1101001000111000  sw	r0, r7
  563=>x"063F",	-- 0000011000111111  dec	r7, r7
  564=>x"D239",	-- 1101001000111001  sw	r1, r7
  565=>x"FFF2",	-- 1111111111110010  liw	r2, font_map
  566=>x"12C0",	-- 0001001011000000  
  567=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  568=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  569=>x"C043",	-- 1100000001000011  li	r3, 8
  570=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  571=>x"0299",	-- 0000001010011001  
  572=>x"D039",	-- 1101000000111001  lw	r1, r7
  573=>x"043F",	-- 0000010000111111  inc	r7, r7
  574=>x"D038",	-- 1101000000111000  lw	r0, r7
  575=>x"043F",	-- 0000010000111111  inc	r7, r7
  576=>x"0400",	-- 0000010000000000  inc	r0, r0
  577=>x"D03E",	-- 1101000000111110  lw	r6, r7
  578=>x"043F",	-- 0000010000111111  inc	r7, r7
  579=>x"E383",	-- 1110001110000011  ba	-, r6
  580=>x"063F",	-- 0000011000111111  dec	r7, r7
  581=>x"D23E",	-- 1101001000111110  sw	r6, r7
  582=>x"FFF4",	-- 1111111111110100  liw	r4, 10000
  583=>x"2710",	-- 0010011100010000  
  584=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  585=>x"0257",	-- 0000001001010111  
  586=>x"FFF4",	-- 1111111111110100  liw	r4, 1000
  587=>x"03E8",	-- 0000001111101000  
  588=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  589=>x"0257",	-- 0000001001010111  
  590=>x"C324",	-- 1100001100100100  li	r4, 100
  591=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  592=>x"0257",	-- 0000001001010111  
  593=>x"C054",	-- 1100000001010100  li	r4, 10
  594=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  595=>x"0257",	-- 0000001001010111  
  596=>x"D03E",	-- 1101000000111110  lw	r6, r7
  597=>x"043F",	-- 0000010000111111  inc	r7, r7
  598=>x"C00C",	-- 1100000000001100  li	r4, 1
  599=>x"C17B",	-- 1100000101111011  li	r3, 0x2F
  600=>x"041B",	-- 0000010000011011  inc	r3, r3
  601=>x"0B12",	-- 0000101100010010  sub	r2, r2, r4
  602=>x"BF91",	-- 1011111110010001  brige	r2, printnum.loop
  603=>x"0912",	-- 0000100100010010  add	r2, r2, r4
  604=>x"063F",	-- 0000011000111111  dec	r7, r7
  605=>x"D23E",	-- 1101001000111110  sw	r6, r7
  606=>x"063F",	-- 0000011000111111  dec	r7, r7
  607=>x"D23A",	-- 1101001000111010  sw	r2, r7
  608=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  609=>x"022F",	-- 0000001000101111  
  610=>x"D03A",	-- 1101000000111010  lw	r2, r7
  611=>x"043F",	-- 0000010000111111  inc	r7, r7
  612=>x"D03E",	-- 1101000000111110  lw	r6, r7
  613=>x"043F",	-- 0000010000111111  inc	r7, r7
  614=>x"E383",	-- 1110001110000011  ba	-, r6
  615=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  616=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  617=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  618=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  619=>x"C0A0",	-- 1100000010100000  li	r0, 20
  620=>x"D011",	-- 1101000000010001  lw	r1, r2
  621=>x"D221",	-- 1101001000100001  sw	r1, r4
  622=>x"0412",	-- 0000010000010010  inc	r2, r2
  623=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  624=>x"061B",	-- 0000011000011011  dec	r3, r3
  625=>x"BEDC",	-- 1011111011011100  brine	r3, put_sprite_16_aligned.loop
  626=>x"E383",	-- 1110001110000011  ba	-, r6
  627=>x"C07D",	-- 1100000001111101  li	r5, 15
  628=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  629=>x"6600",	-- 0110011000000000  shr	r0, r0, 3
  630=>x"BC68",	-- 1011110001101000  brieq	r5, put_sprite_16_aligned
  631=>x"062D",	-- 0000011000101101  dec	r5, r5
  632=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  633=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  634=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  635=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  636=>x"063F",	-- 0000011000111111  dec	r7, r7
  637=>x"D23B",	-- 1101001000111011  sw	r3, r7
  638=>x"D011",	-- 1101000000010001  lw	r1, r2
  639=>x"CFF8",	-- 1100111111111000  li	r0, -1
  640=>x"3D40",	-- 0011110101000000  rsr	r0, r0, r5
  641=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  642=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  643=>x"D023",	-- 1101000000100011  lw	r3, r4
  644=>x"2600",	-- 0010011000000000  not	r0, r0
  645=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  646=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  647=>x"D221",	-- 1101001000100001  sw	r1, r4
  648=>x"0424",	-- 0000010000100100  inc	r4, r4
  649=>x"D011",	-- 1101000000010001  lw	r1, r2
  650=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  651=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  652=>x"D023",	-- 1101000000100011  lw	r3, r4
  653=>x"2600",	-- 0010011000000000  not	r0, r0
  654=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  655=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  656=>x"D221",	-- 1101001000100001  sw	r1, r4
  657=>x"0412",	-- 0000010000010010  inc	r2, r2
  658=>x"C098",	-- 1100000010011000  li	r0, 19
  659=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  660=>x"D03B",	-- 1101000000111011  lw	r3, r7
  661=>x"043F",	-- 0000010000111111  inc	r7, r7
  662=>x"061B",	-- 0000011000011011  dec	r3, r3
  663=>x"B95C",	-- 1011100101011100  brine	r3, put_sprite_16.loop
  664=>x"E383",	-- 1110001110000011  ba	-, r6
  665=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  666=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  667=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  668=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  669=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  670=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  671=>x"C0A5",	-- 1100000010100101  li	r5, 20
  672=>x"8404",	-- 1000010000000100  brine	r0, put_sprite_8_aligned.loop1
  673=>x"D010",	-- 1101000000010000  lw	r0, r2
  674=>x"D021",	-- 1101000000100001  lw	r1, r4
  675=>x"1A41",	-- 0001101001000001  mixhl	r1, r0, r1
  676=>x"D221",	-- 1101001000100001  sw	r1, r4
  677=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  678=>x"061B",	-- 0000011000011011  dec	r3, r3
  679=>x"E398",	-- 1110001110011000  baeq	r3, r6
  680=>x"D021",	-- 1101000000100001  lw	r1, r4
  681=>x"1E41",	-- 0001111001000001  mixll	r1, r0, r1
  682=>x"D221",	-- 1101001000100001  sw	r1, r4
  683=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  684=>x"0412",	-- 0000010000010010  inc	r2, r2
  685=>x"061B",	-- 0000011000011011  dec	r3, r3
  686=>x"E398",	-- 1110001110011000  baeq	r3, r6
  687=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop0
  688=>x"D010",	-- 1101000000010000  lw	r0, r2
  689=>x"D021",	-- 1101000000100001  lw	r1, r4
  690=>x"1809",	-- 0001100000001001  mixhh	r1, r1, r0
  691=>x"D221",	-- 1101001000100001  sw	r1, r4
  692=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  693=>x"061B",	-- 0000011000011011  dec	r3, r3
  694=>x"E398",	-- 1110001110011000  baeq	r3, r6
  695=>x"D021",	-- 1101000000100001  lw	r1, r4
  696=>x"1A09",	-- 0001101000001001  mixhl	r1, r1, r0
  697=>x"D221",	-- 1101001000100001  sw	r1, r4
  698=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  699=>x"0412",	-- 0000010000010010  inc	r2, r2
  700=>x"061B",	-- 0000011000011011  dec	r3, r3
  701=>x"E398",	-- 1110001110011000  baeq	r3, r6
  702=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop1
  703=>x"C03D",	-- 1100000000111101  li	r5, 7
  704=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  705=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  706=>x"B5E8",	-- 1011010111101000  brieq	r5, put_sprite_8_aligned
  707=>x"062D",	-- 0000011000101101  dec	r5, r5
  708=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  709=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  710=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  711=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  712=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  713=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  714=>x"8A04",	-- 1000101000000100  brine	r0, put_sprite_8.loop1
  715=>x"D010",	-- 1101000000010000  lw	r0, r2
  716=>x"063F",	-- 0000011000111111  dec	r7, r7
  717=>x"D23A",	-- 1101001000111010  sw	r2, r7
  718=>x"C802",	-- 1100100000000010  li	r2, 0x100
  719=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  720=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  721=>x"D021",	-- 1101000000100001  lw	r1, r4
  722=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  723=>x"2612",	-- 0010011000010010  not	r2, r2
  724=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  725=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  726=>x"D221",	-- 1101001000100001  sw	r1, r4
  727=>x"C0A1",	-- 1100000010100001  li	r1, 20
  728=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  729=>x"D03A",	-- 1101000000111010  lw	r2, r7
  730=>x"043F",	-- 0000010000111111  inc	r7, r7
  731=>x"061B",	-- 0000011000011011  dec	r3, r3
  732=>x"E398",	-- 1110001110011000  baeq	r3, r6
  733=>x"D010",	-- 1101000000010000  lw	r0, r2
  734=>x"063F",	-- 0000011000111111  dec	r7, r7
  735=>x"D23A",	-- 1101001000111010  sw	r2, r7
  736=>x"1E00",	-- 0001111000000000  mixll	r0, r0, r0
  737=>x"C802",	-- 1100100000000010  li	r2, 0x100
  738=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  739=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  740=>x"D021",	-- 1101000000100001  lw	r1, r4
  741=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  742=>x"2612",	-- 0010011000010010  not	r2, r2
  743=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  744=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  745=>x"D221",	-- 1101001000100001  sw	r1, r4
  746=>x"C0A1",	-- 1100000010100001  li	r1, 20
  747=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  748=>x"D03A",	-- 1101000000111010  lw	r2, r7
  749=>x"043F",	-- 0000010000111111  inc	r7, r7
  750=>x"0412",	-- 0000010000010010  inc	r2, r2
  751=>x"061B",	-- 0000011000011011  dec	r3, r3
  752=>x"E398",	-- 1110001110011000  baeq	r3, r6
  753=>x"B683",	-- 1011011010000011  bri	-, put_sprite_8.loop0
  754=>x"D010",	-- 1101000000010000  lw	r0, r2
  755=>x"063F",	-- 0000011000111111  dec	r7, r7
  756=>x"D23A",	-- 1101001000111010  sw	r2, r7
  757=>x"063F",	-- 0000011000111111  dec	r7, r7
  758=>x"D23B",	-- 1101001000111011  sw	r3, r7
  759=>x"C802",	-- 1100100000000010  li	r2, 0x100
  760=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  761=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  762=>x"2080",	-- 0010000010000000  and	r0, r0, r2
  763=>x"D021",	-- 1101000000100001  lw	r1, r4
  764=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
  765=>x"261B",	-- 0010011000011011  not	r3, r3
  766=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  767=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
  768=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  769=>x"D221",	-- 1101001000100001  sw	r1, r4
  770=>x"0424",	-- 0000010000100100  inc	r4, r4
  771=>x"D021",	-- 1101000000100001  lw	r1, r4
  772=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  773=>x"261B",	-- 0010011000011011  not	r3, r3
  774=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  775=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
  776=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  777=>x"D221",	-- 1101001000100001  sw	r1, r4
  778=>x"C099",	-- 1100000010011001  li	r1, 19
  779=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  780=>x"D03B",	-- 1101000000111011  lw	r3, r7
  781=>x"043F",	-- 0000010000111111  inc	r7, r7
  782=>x"D03A",	-- 1101000000111010  lw	r2, r7
  783=>x"043F",	-- 0000010000111111  inc	r7, r7
  784=>x"061B",	-- 0000011000011011  dec	r3, r3
  785=>x"E398",	-- 1110001110011000  baeq	r3, r6
  786=>x"D010",	-- 1101000000010000  lw	r0, r2
  787=>x"4E00",	-- 0100111000000000  shl	r0, r0, 7
  788=>x"063F",	-- 0000011000111111  dec	r7, r7
  789=>x"D23A",	-- 1101001000111010  sw	r2, r7
  790=>x"063F",	-- 0000011000111111  dec	r7, r7
  791=>x"D23B",	-- 1101001000111011  sw	r3, r7
  792=>x"C802",	-- 1100100000000010  li	r2, 0x100
  793=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  794=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  795=>x"2080",	-- 0010000010000000  and	r0, r0, r2
  796=>x"D021",	-- 1101000000100001  lw	r1, r4
  797=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
  798=>x"261B",	-- 0010011000011011  not	r3, r3
  799=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  800=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
  801=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  802=>x"D221",	-- 1101001000100001  sw	r1, r4
  803=>x"0424",	-- 0000010000100100  inc	r4, r4
  804=>x"D021",	-- 1101000000100001  lw	r1, r4
  805=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  806=>x"261B",	-- 0010011000011011  not	r3, r3
  807=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  808=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
  809=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  810=>x"D221",	-- 1101001000100001  sw	r1, r4
  811=>x"C099",	-- 1100000010011001  li	r1, 19
  812=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  813=>x"D03B",	-- 1101000000111011  lw	r3, r7
  814=>x"043F",	-- 0000010000111111  inc	r7, r7
  815=>x"D03A",	-- 1101000000111010  lw	r2, r7
  816=>x"043F",	-- 0000010000111111  inc	r7, r7
  817=>x"0412",	-- 0000010000010010  inc	r2, r2
  818=>x"061B",	-- 0000011000011011  dec	r3, r3
  819=>x"E398",	-- 1110001110011000  baeq	r3, r6
  820=>x"AF83",	-- 1010111110000011  bri	-, put_sprite_8.loop1
    others => x"0000"
    );
begin
  process(CLK)
  begin
    if (CLK'event AND CLK='1') then
      D <= m(to_integer(unsigned(AD)));
    end if;
  end process;
end Behavioral;
