----------------------------------------------------------------------------------
--
-- File retrieved, on 07/02/2010, from :
-- http://sebastien-viardot.imag.fr/Enseignements/Archi1A2s/sources/ROMPROG.vhd
--
-- Slightly altered to get rid of vendor-specific packages and adjust formatting
--
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROMPROG is
  Port ( AD : in  STD_LOGIC_VECTOR (12 downto 0);
         D : out  STD_LOGIC_VECTOR (15 downto 0);
         CLK : in STD_LOGIC);
end ROMPROG;

architecture Behavioral of ROMPROG is
  constant low_address: natural := 0;
  constant high_address: natural := 8192;
  subtype octet is std_logic_vector( 15 downto 0 );
  type zone_memoire is
    array (natural range low_address to high_address-1) of octet;
  constant m: zone_memoire:= (
0=>x"25FF",     -- 0010010111111111  xor        r7, r7, r7
1=>x"F8C0",     -- 1111100011000000  bai        -, os_init
2=>x"0100",     -- 0000000100000000  

16=>x"FFF0",    -- 1111111111110000  liw        r0, IRQ_ack
17=>x"2002",    -- 0010000000000010  
18=>x"CFF9",    -- 1100111111111001  li r1, -1
19=>x"D201",    -- 1101001000000001  sw r1, r0
20=>x"261B",    -- 0010011000011011  not r3, r3
21=>x"D6C0",    -- 1101011011000000  out        r3
22=>x"FFFE",    -- 1111111111111110  reti

256=>x"FFF0",   -- 1111111111110000  liw        r0, IRQ_mask
257=>x"2000",   -- 0010000000000000  
258=>x"C009",   -- 1100000000001001  li r1, 1
259=>x"D201",   -- 1101001000000001  sw r1, r0
260=>x"0400",   -- 0000010000000000  inc        r0, r0
261=>x"CFF9",   -- 1100111111111001  li r1, -1
262=>x"D201",   -- 1101001000000001  sw r1, r0
263=>x"C03A",   -- 1100000000111010  li r2, 7
264=>x"0880",   -- 0000100010000000  add        r0, r0, r2
265=>x"C0F2",   -- 1100000011110010  li r2, 0x1E
266=>x"D202",   -- 1101001000000010  sw r2, r0
267=>x"0400",   -- 0000010000000000  inc        r0, r0
268=>x"C012",   -- 1100000000010010  li r2, 2
269=>x"D202",   -- 1101001000000010  sw r2, r0

270=>x"FFF0",   -- 1111111111110000  liw        r0, 0x8421
271=>x"8421",   -- 1000010000100001  
272=>x"FFF1",   -- 1111111111110001  liw        r1, 0x1234
273=>x"1234",   -- 0001001000110100  
274=>x"E408",   -- 1110010000001000  exw        r0, r1
275=>x"E408",   -- 1110010000001000  exw        r0, r1
276=>x"1842",   -- 0001100001000010  mixhh      r2, r0, r1
277=>x"1A43",   -- 0001101001000011  mixhl      r3, r0, r1
278=>x"1C44",   -- 0001110001000100  mixlh      r4, r0, r1
279=>x"1E45",   -- 0001111001000101  mixll      r5, r0, r1

280=>x"C000",   -- 1100000000000000  li r0, 0
281=>x"C001",   -- 1100000000000001  li r1, 0
282=>x"FFF2",   -- 1111111111110010  liw        r2, hello_str
283=>x"16C0",   -- 0001011011000000  
284=>x"FAC6",   -- 1111101011000110  bail       -, r6, puts
285=>x"014F",   -- 0000000101001111  

286=>x"C750",   -- 1100011101010000  li r0, 234
287=>x"C1C2",   -- 1100000111000010  li r2, 56
288=>x"FAC6",   -- 1111101011000110  bail       -, r6, div_16_16
289=>x"0138",   -- 0000000100111000  

290=>x"C448",   -- 1100010001001000  li r0, 137
291=>x"C472",   -- 1100010001110010  li r2, 142
292=>x"FAC6",   -- 1111101011000110  bail       -, r6, mult_16_16
293=>x"012C",   -- 0000000100101100  

294=>x"C03A",   -- 1100000000111010  li r2, 7
295=>x"FAC6",   -- 1111101011000110  bail       -, r6, fact_16
296=>x"0143",   -- 0000000101000011  

297=>x"C079",   -- 1100000001111001  li r1, 15
298=>x"2008",   -- 0010000000001000  and        r0, r1, r0
299=>x"BB83",   -- 1011101110000011  bri        -, test.puts + 1

300=>x"2449",   -- 0010010001001001  xor        r1, r1, r1
301=>x"2524",   -- 0010010100100100  xor        r4, r4, r4
302=>x"C085",   -- 1100000010000101  li r5, 16
303=>x"0849",   -- 0000100001001001  add        r1, r1, r1
304=>x"0C00",   -- 0000110000000000  adc        r0, r0, r0
305=>x"0EDB",   -- 0000111011011011  sbc        r3, r3, r3
306=>x"209B",   -- 0010000010011011  and        r3, r3, r2
307=>x"08C9",   -- 0000100011001001  add        r1, r1, r3
308=>x"0D00",   -- 0000110100000000  adc        r0, r0, r4
309=>x"062D",   -- 0000011000101101  dec        r5, r5
310=>x"BE6C",   -- 1011111001101100  brine      r5, mult_16_16.loop
311=>x"E383",   -- 1110001110000011  ba -, r6

312=>x"2449",   -- 0010010001001001  xor        r1, r1, r1
313=>x"C084",   -- 1100000010000100  li r4, 16
314=>x"0800",   -- 0000100000000000  add        r0, r0, r0
315=>x"0C49",   -- 0000110001001001  adc        r1, r1, r1
316=>x"0A8B",   -- 0000101010001011  sub        r3, r1, r2
317=>x"80DD",   -- 1000000011011101  brilt      r3, div_16_16.skip
318=>x"0A89",   -- 0000101010001001  sub        r1, r1, r2
319=>x"0400",   -- 0000010000000000  inc        r0, r0
320=>x"0624",   -- 0000011000100100  dec        r4, r4
321=>x"BE64",   -- 1011111001100100  brine      r4, div_16_16.loop
322=>x"E383",   -- 1110001110000011  ba -, r6

323=>x"2400",   -- 0010010000000000  xor        r0, r0, r0
324=>x"2449",   -- 0010010001001001  xor        r1, r1, r1
325=>x"8250",   -- 1000001001010000  brieq      r2, fact_16.end
326=>x"0409",   -- 0000010000001001  inc        r1, r1
327=>x"1008",   -- 0001000000001000  mova       r0, r1
328=>x"FAC6",   -- 1111101011000110  bail       -, r6, mult_16_16
329=>x"012C",   -- 0000000100101100  
330=>x"8104",   -- 1000000100000100  brine      r0, fact_16.overflow
331=>x"012C",   -- 0000000100101100  
332=>x"0612",   -- 0000011000010010  dec        r2, r2
333=>x"BE94",   -- 1011111010010100  brine      r2, fact_16.loop
334=>x"E383",   -- 1110001110000011  ba -, r6

335=>x"D013",   -- 1101000000010011  lw r3, r2
336=>x"6E1B",   -- 0110111000011011  shr        r3, r3, 7
337=>x"E398",   -- 1110001110011000  baeq       r3, r6
338=>x"063F",   -- 0000011000111111  dec        r7, r7
339=>x"D23E",   -- 1101001000111110  sw r6, r7
340=>x"063F",   -- 0000011000111111  dec        r7, r7
341=>x"D238",   -- 1101001000111000  sw r0, r7
342=>x"063F",   -- 0000011000111111  dec        r7, r7
343=>x"D239",   -- 1101001000111001  sw r1, r7
344=>x"063F",   -- 0000011000111111  dec        r7, r7
345=>x"D23A",   -- 1101001000111010  sw r2, r7
346=>x"FFF4",   -- 1111111111110100  liw        r4, font_map
347=>x"12C0",   -- 0001001011000000  
348=>x"091A",   -- 0000100100011010  add        r2, r3, r4
349=>x"C043",   -- 1100000001000011  li r3, 8
350=>x"FAC6",   -- 1111101011000110  bail       -, r6, put_sprite_8_aligned
351=>x"018D",   -- 0000000110001101  
352=>x"D03A",   -- 1101000000111010  lw r2, r7
353=>x"043F",   -- 0000010000111111  inc        r7, r7
354=>x"D039",   -- 1101000000111001  lw r1, r7
355=>x"043F",   -- 0000010000111111  inc        r7, r7
356=>x"D038",   -- 1101000000111000  lw r0, r7
357=>x"043F",   -- 0000010000111111  inc        r7, r7
358=>x"0400",   -- 0000010000000000  inc        r0, r0
359=>x"D013",   -- 1101000000010011  lw r3, r2
360=>x"4E1B",   -- 0100111000011011  shl        r3, r3, 7
361=>x"6E1B",   -- 0110111000011011  shr        r3, r3, 7
362=>x"E398",   -- 1110001110011000  baeq       r3, r6
363=>x"063F",   -- 0000011000111111  dec        r7, r7
364=>x"D238",   -- 1101001000111000  sw r0, r7
365=>x"063F",   -- 0000011000111111  dec        r7, r7
366=>x"D239",   -- 1101001000111001  sw r1, r7
367=>x"063F",   -- 0000011000111111  dec        r7, r7
368=>x"D23A",   -- 1101001000111010  sw r2, r7
369=>x"FFF4",   -- 1111111111110100  liw        r4, font_map
370=>x"12C0",   -- 0001001011000000  
371=>x"091A",   -- 0000100100011010  add        r2, r3, r4
372=>x"C043",   -- 1100000001000011  li r3, 8
373=>x"FAC6",   -- 1111101011000110  bail       -, r6, put_sprite_8_aligned
374=>x"018D",   -- 0000000110001101  
375=>x"D03A",   -- 1101000000111010  lw r2, r7
376=>x"043F",   -- 0000010000111111  inc        r7, r7
377=>x"D039",   -- 1101000000111001  lw r1, r7
378=>x"043F",   -- 0000010000111111  inc        r7, r7
379=>x"D038",   -- 1101000000111000  lw r0, r7
380=>x"043F",   -- 0000010000111111  inc        r7, r7
381=>x"0400",   -- 0000010000000000  inc        r0, r0
382=>x"D03E",   -- 1101000000111110  lw r6, r7
383=>x"043F",   -- 0000010000111111  inc        r7, r7
384=>x"0412",   -- 0000010000010010  inc        r2, r2
385=>x"B383",   -- 1011001110000011  bri        -, puts.loop

386=>x"460C",   -- 0100011000001100  shl r4, r1, 3
387=>x"4209",   -- 0100001000001001  shl        r1, r1, 1
388=>x"0864",   -- 0000100001100100  add        r4, r4, r1
389=>x"0824",   -- 0000100000100100  add        r4, r4, r0
390=>x"D011",   -- 1101000000010001  lw r1, r2
391=>x"D221",   -- 1101001000100001  sw r1, r4
392=>x"0412",   -- 0000010000010010  inc        r2, r2
393=>x"0424",   -- 0000010000100100  inc        r4, r4
394=>x"061B",   -- 0000011000011011  dec        r3, r3
395=>x"BEDC",   -- 1011111011011100  brine      r3, put_sprite_16_aligned.loop
396=>x"E383",   -- 1110001110000011  ba -, r6

397=>x"460C",   -- 0100011000001100  shl r4, r1, 3
398=>x"4209",   -- 0100001000001001  shl        r1, r1, 1
399=>x"0864",   -- 0000100001100100  add        r4, r4, r1
400=>x"4001",   -- 0100000000000001  shl        r1, r0, 0
401=>x"0E00",   -- 0000111000000000  sbc        r0, r0, r0
402=>x"0864",   -- 0000100001100100  add        r4, r4, r1
403=>x"C0A5",   -- 1100000010100101  li r5, 20
404=>x"83C4",   -- 1000001111000100  brine      r0, put_sprite_8_aligned.loop1
405=>x"D010",   -- 1101000000010000  lw r0, r2
406=>x"D021",   -- 1101000000100001  lw r1, r4
407=>x"1A41",   -- 0001101001000001  mixhl      r1, r0, r1
408=>x"D221",   -- 1101001000100001  sw r1, r4
409=>x"061B",   -- 0000011000011011  dec        r3, r3
410=>x"8218",   -- 1000001000011000  brieq      r3, put_sprite_8_aligned.end
411=>x"0964",   -- 0000100101100100  add        r4, r4, r5
412=>x"D021",   -- 1101000000100001  lw r1, r4
413=>x"1E41",   -- 0001111001000001  mixll      r1, r0, r1
414=>x"D221",   -- 1101001000100001  sw r1, r4
415=>x"0412",   -- 0000010000010010  inc        r2, r2
416=>x"061B",   -- 0000011000011011  dec        r3, r3
417=>x"BD1C",   -- 1011110100011100  brine      r3, put_sprite_8_aligned.loop0
418=>x"E383",   -- 1110001110000011  ba -, r6
419=>x"D010",   -- 1101000000010000  lw r0, r2
420=>x"D021",   -- 1101000000100001  lw r1, r4
421=>x"1809",   -- 0001100000001001  mixhh      r1, r1, r0
422=>x"D221",   -- 1101001000100001  sw r1, r4
423=>x"061B",   -- 0000011000011011  dec        r3, r3
424=>x"BE98",   -- 1011111010011000  brieq      r3, put_sprite_8_aligned.end
425=>x"0964",   -- 0000100101100100  add        r4, r4, r5
426=>x"D021",   -- 1101000000100001  lw r1, r4
427=>x"1A09",   -- 0001101000001001  mixhl      r1, r1, r0
428=>x"D221",   -- 1101001000100001  sw r1, r4
429=>x"0412",   -- 0000010000010010  inc        r2, r2
430=>x"061B",   -- 0000011000011011  dec        r3, r3
431=>x"BD1C",   -- 1011110100011100  brine      r3, put_sprite_8_aligned.loop1
432=>x"E383",   -- 1110001110000011  ba -, r6

--     0=>X"D400", -- IN R0
--     1=>X"D600", -- OUT R0
--     2=>X"8043", -- bri r0, 1
--     3=>X"D400", -- IN R0
--     4=>X"D600", -- OUT R0
--     5=>X"FFFF", -- RESET
    others => x"0000"
    );
begin
  process(CLK)
  begin
    if (CLK'event AND CLK='1') then
      D <= m(to_integer(unsigned(AD)));
    end if;
  end process;
end Behavioral;
