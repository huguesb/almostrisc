----------------------------------------------------------------------------------
--
-- File retrieved, on 07/02/2010, from :
-- http://sebastien-viardot.imag.fr/Enseignements/Archi1A2s/sources/ROMPROG.vhd
--
-- Slightly altered to get rid of vendor-specific packages and adjust formatting
-- Now auto-filled by asrom script
--
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROMPROG is
  Port ( AD : in  STD_LOGIC_VECTOR (12 downto 0);
         D : out  STD_LOGIC_VECTOR (15 downto 0);
         CLK : in STD_LOGIC);
end ROMPROG;

architecture Behavioral of ROMPROG is
  constant low_address: natural := 0;
  constant high_address: natural := 8192;
  subtype octet is std_logic_vector( 15 downto 0 );
  type zone_memoire is
    array (natural range low_address to high_address-1) of octet;
  constant m: zone_memoire:= (
    0=>x"FFF7",	-- 1111111111110111  liw	r7, IRQ_mask
    1=>x"2000",	-- 0010000000000000  
    2=>x"F8C0",	-- 1111100011000000  bai	-, os_init
    3=>x"0100",	-- 0000000100000000  
   16=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_ack
   17=>x"2002",	-- 0010000000000010  
   18=>x"D001",	-- 1101000000000001  lw	r1, r0
   19=>x"F54A",	-- 1111010101001010  bspl	r2, r1, 5
   20=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_error
   21=>x"0050",	-- 0000000001010000  
   22=>x"F4CA",	-- 1111010011001010  bspl	r2, r1, 3
   23=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_kbd
   24=>x"0060",	-- 0000000001100000  
   25=>x"F40A",	-- 1111010000001010  bspl	r2, r1, 0
   26=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_tmr
   27=>x"0040",	-- 0000000001000000  
   28=>x"D201",	-- 1101001000000001  sw	r1, r0
   29=>x"FFFE",	-- 1111111111111110  reti
   64=>x"263F",	-- 0010011000111111  not r7, r7
   65=>x"D7C0",	-- 1101011111000000  out	r7
   66=>x"E383",	-- 1110001110000011  ba	-, r6
   80=>x"25FF",	-- 0010010111111111  xor	r7, r7, r7
   81=>x"D7C0",	-- 1101011111000000  out	r7
   82=>x"E383",	-- 1110001110000011  ba	-, r6
   96=>x"FFF2",	-- 1111111111110010  liw	r2, PS2_rx
   97=>x"2004",	-- 0010000000000100  
   98=>x"D012",	-- 1101000000010010  lw	r2, r2
   99=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map + 8
  100=>x"16C8",	-- 0001011011001000  
  101=>x"D01B",	-- 1101000000011011  lw	r3, r3
  102=>x"1EBF",	-- 0001111010111111  mixll	r7, r7, r2
  103=>x"C784",	-- 1100011110000100  li	r4, 0xF0
  104=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  105=>x"8B20",	-- 1000101100100000  brieq	r4, int_kbd.release
  106=>x"C704",	-- 1100011100000100  li	r4, 0xE0
  107=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  108=>x"88E0",	-- 1000100011100000  brieq	r4, int_kbd.extended
  109=>x"FFF5",	-- 1111111111110101  liw	r5, paper_keys - 1
  110=>x"16CF",	-- 0001011011001111  
  111=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  112=>x"80E0",	-- 1000000011100000  brieq	r4, $+3
  113=>x"FFF5",	-- 1111111111110101  liw	r5, paper_keys + 11 - 1
  114=>x"16DA",	-- 0001011011011010  
  115=>x"042D",	-- 0000010000101101  inc	r5, r5
  116=>x"D02C",	-- 1101000000101100  lw	r4, r5
  117=>x"8560",	-- 1000010101100000  brieq	r4, scan_code_mismatch
  118=>x"6E24",	-- 0110111000100100  shr	r4, r4, 7
  119=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  120=>x"BEE4",	-- 1011111011100100  brine	r4, scan_code_loop
  121=>x"D02A",	-- 1101000000101010  lw	r2, r5
  122=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  123=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  124=>x"741B",	-- 0111010000011011  shr	r3, r3, 10
  125=>x"C00D",	-- 1100000000001101  li	r5, 1
  126=>x"0612",	-- 0000011000010010  dec	r2, r2
  127=>x"3AAA",	-- 0011101010101010  rrl	r2, r5, r2
  128=>x"FFF5",	-- 1111111111110101  liw	r5, key_press_map
  129=>x"16C0",	-- 0001011011000000  
  130=>x"08ED",	-- 0000100011101101  add	r5, r5, r3
  131=>x"D02B",	-- 1101000000101011  lw	r3, r5
  132=>x"80E4",	-- 1000000011100100  brine	r4, scan_code_release
  133=>x"229B",	-- 0010001010011011  or	r3, r3, r2
  134=>x"80C3",	-- 1000000011000011  bri	-, scan_code_notify
  135=>x"2612",	-- 0010011000010010  not	r2, r2
  136=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  137=>x"D22B",	-- 1101001000101011  sw	r3, r5
  138=>x"C003",	-- 1100000000000011  li	r3, 0
  139=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  140=>x"16C8",	-- 0001011011001000  
  141=>x"D223",	-- 1101001000100011  sw	r3, r4
  142=>x"E383",	-- 1110001110000011  ba	-, r6
  143=>x"C014",	-- 1100000000010100  li	r4, 2
  144=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  145=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  146=>x"16C8",	-- 0001011011001000  
  147=>x"D223",	-- 1101001000100011  sw	r3, r4
  148=>x"E383",	-- 1110001110000011  ba	-, r6
  149=>x"C00C",	-- 1100000000001100  li	r4, 1
  150=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  151=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  152=>x"16C8",	-- 0001011011001000  
  153=>x"D223",	-- 1101001000100011  sw	r3, r4
  154=>x"E383",	-- 1110001110000011  ba	-, r6
  256=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_mask
  257=>x"2000",	-- 0010000000000000  
  258=>x"C0C9",	-- 1100000011001001  li	r1, 0x19
  259=>x"D201",	-- 1101001000000001  sw	r1, r0
  260=>x"0400",	-- 0000010000000000  inc	r0, r0
  261=>x"CFF9",	-- 1100111111111001  li	r1, -1
  262=>x"D201",	-- 1101001000000001  sw	r1, r0
  263=>x"C03A",	-- 1100000000111010  li	r2, 7
  264=>x"0880",	-- 0000100010000000  add	r0, r0, r2
  265=>x"C0EA",	-- 1100000011101010  li	r2, 0x1D
  266=>x"D202",	-- 1101001000000010  sw	r2, r0
  267=>x"0400",	-- 0000010000000000  inc	r0, r0
  268=>x"C07A",	-- 1100000001111010  li	r2, 15
  269=>x"D202",	-- 1101001000000010  sw	r2, r0
  270=>x"0400",	-- 0000010000000000  inc	r0, r0
  271=>x"C0DA",	-- 1100000011011010  li	r2, 0x1B
  272=>x"D202",	-- 1101001000000010  sw	r2, r0
  273=>x"0400",	-- 0000010000000000  inc	r0, r0
  274=>x"FFF2",	-- 1111111111110010  liw	r2, 817
  275=>x"0331",	-- 0000001100110001  
  276=>x"D202",	-- 1101001000000010  sw	r2, r0
  277=>x"FFF0",	-- 1111111111110000  liw	r0, key_press_map
  278=>x"16C0",	-- 0001011011000000  
  279=>x"C001",	-- 1100000000000001  li	r1, 0
  280=>x"C042",	-- 1100000001000010  li	r2, 8
  281=>x"D201",	-- 1101001000000001  sw	r1, r0
  282=>x"0400",	-- 0000010000000000  inc	r0, r0
  283=>x"0612",	-- 0000011000010010  dec	r2, r2
  284=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  285=>x"C0F3",	-- 1100000011110011  li	r3, 30
  286=>x"CFFA",	-- 1100111111111010  li	r2, -1
  287=>x"D21A",	-- 1101001000011010  sw	r2, r3
  288=>x"8083",	-- 1000000010000011  bri	-, PaperGameStart
  289=>x"8003",	-- 1000000000000011  bri	-, PaperMenuLoop
  290=>x"FFF0",	-- 1111111111110000  liw	r0, paper_dir
  291=>x"179C",	-- 0001011110011100  
  292=>x"C001",	-- 1100000000000001  li	r1, 0
  293=>x"D201",	-- 1101001000000001  sw	r1, r0
  294=>x"0400",	-- 0000010000000000  inc	r0, r0
  295=>x"FFF1",	-- 1111111111110001  liw	r1, 152 * 8
  296=>x"04C0",	-- 0000010011000000  
  297=>x"D201",	-- 1101001000000001  sw	r1, r0
  298=>x"0400",	-- 0000010000000000  inc	r0, r0
  299=>x"C001",	-- 1100000000000001  li	r1, 0
  300=>x"D201",	-- 1101001000000001  sw	r1, r0
  301=>x"0400",	-- 0000010000000000  inc	r0, r0
  302=>x"FFF1",	-- 1111111111110001  liw	r1, 128 * 8
  303=>x"0400",	-- 0000010000000000  
  304=>x"D201",	-- 1101001000000001  sw	r1, r0
  305=>x"0400",	-- 0000010000000000  inc	r0, r0
  306=>x"C001",	-- 1100000000000001  li	r1, 0
  307=>x"D201",	-- 1101001000000001  sw	r1, r0
  308=>x"0400",	-- 0000010000000000  inc	r0, r0
  309=>x"C029",	-- 1100000000101001  li	r1, 5
  310=>x"D201",	-- 1101001000000001  sw	r1, r0
  311=>x"0400",	-- 0000010000000000  inc	r0, r0
  312=>x"C011",	-- 1100000000010001  li	r1, 2
  313=>x"D201",	-- 1101001000000001  sw	r1, r0
  314=>x"0400",	-- 0000010000000000  inc	r0, r0
  315=>x"FFF0",	-- 1111111111110000  liw	r0, TMR_cur1
  316=>x"200D",	-- 0010000000001101  
  317=>x"D000",	-- 1101000000000000  lw	r0, r0
  318=>x"FAC6",	-- 1111101011000110  bail	-, r6, rand16_init
  319=>x"0221",	-- 0000001000100001  
  320=>x"C000",	-- 1100000000000000  li	r0, 0
  321=>x"CFF9",	-- 1100111111111001  li	r1, -1
  322=>x"C0A2",	-- 1100000010100010  li	r2, 20
  323=>x"D201",	-- 1101001000000001  sw	r1, r0
  324=>x"0400",	-- 0000010000000000  inc	r0, r0
  325=>x"0612",	-- 0000011000010010  dec	r2, r2
  326=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  327=>x"C001",	-- 1100000000000001  li	r1, 0
  328=>x"FFF2",	-- 1111111111110010  liw	r2, 18*20
  329=>x"0168",	-- 0000000101101000  
  330=>x"D201",	-- 1101001000000001  sw	r1, r0
  331=>x"0400",	-- 0000010000000000  inc	r0, r0
  332=>x"0612",	-- 0000011000010010  dec	r2, r2
  333=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  334=>x"CFF9",	-- 1100111111111001  li	r1, -1
  335=>x"C0A2",	-- 1100000010100010  li	r2, 20
  336=>x"D201",	-- 1101001000000001  sw	r1, r0
  337=>x"0400",	-- 0000010000000000  inc	r0, r0
  338=>x"0612",	-- 0000011000010010  dec	r2, r2
  339=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  340=>x"C020",	-- 1100000000100000  li	r0, 4
  341=>x"C029",	-- 1100000000101001  li	r1, 5
  342=>x"FFF2",	-- 1111111111110010  liw	r2, paper_title
  343=>x"17A4",	-- 0001011110100100  
  344=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  345=>x"0267",	-- 0000001001100111  
  346=>x"C778",	-- 1100011101111000  li	r0, 239
  347=>x"C009",	-- 1100000000001001  li	r1, 1
  348=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud
  349=>x"1780",	-- 0001011110000000  
  350=>x"C043",	-- 1100000001000011  li	r3, 8
  351=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  352=>x"0356",	-- 0000001101010110  
  353=>x"C0F8",	-- 1100000011111000  li	r0, 31
  354=>x"C009",	-- 1100000000001001  li	r1, 1
  355=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed + 1
  356=>x"17A1",	-- 0001011110100001  
  357=>x"D012",	-- 1101000000010010  lw	r2, r2
  358=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum
  359=>x"0296",	-- 0000001010010110  
  360=>x"C120",	-- 1100000100100000  li	r0, 36
  361=>x"C009",	-- 1100000000001001  li	r1, 1
  362=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  363=>x"17AA",	-- 0001011110101010  
  364=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  365=>x"0267",	-- 0000001001100111  
  366=>x"C778",	-- 1100011101111000  li	r0, 239
  367=>x"C051",	-- 1100000001010001  li	r1, 10
  368=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud + 4
  369=>x"1784",	-- 0001011110000100  
  370=>x"C043",	-- 1100000001000011  li	r3, 8
  371=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  372=>x"0356",	-- 0000001101010110  
  373=>x"C0F8",	-- 1100000011111000  li	r0, 31
  374=>x"C051",	-- 1100000001010001  li	r1, 10
  375=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed + 2
  376=>x"17A2",	-- 0001011110100010  
  377=>x"D012",	-- 1101000000010010  lw	r2, r2
  378=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum
  379=>x"0296",	-- 0000001010010110  
  380=>x"C120",	-- 1100000100100000  li	r0, 36
  381=>x"C051",	-- 1100000001010001  li	r1, 10
  382=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  383=>x"17AA",	-- 0001011110101010  
  384=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  385=>x"0267",	-- 0000001001100111  
  386=>x"FFF0",	-- 1111111111110000  liw	r0, 20*20
  387=>x"0190",	-- 0000000110010000  
  388=>x"C001",	-- 1100000000000001  li	r1, 0
  389=>x"FFF2",	-- 1111111111110010  liw	r2, 220*20
  390=>x"1130",	-- 0001000100110000  
  391=>x"D201",	-- 1101001000000001  sw	r1, r0
  392=>x"0400",	-- 0000010000000000  inc	r0, r0
  393=>x"0612",	-- 0000011000010010  dec	r2, r2
  394=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  395=>x"FFF5",	-- 1111111111110101  liw	r5, paper_tilemap
  396=>x"17B0",	-- 0001011110110000  
  397=>x"D02C",	-- 1101000000101100  lw	r4, r5
  398=>x"042D",	-- 0000010000101101  inc	r5, r5
  399=>x"88E0",	-- 1000100011100000  brieq	r4, PaperGameTileSkip
  400=>x"063F",	-- 0000011000111111  dec	r7, r7
  401=>x"D23D",	-- 1101001000111101  sw	r5, r7
  402=>x"FFF3",	-- 1111111111110011  liw	r3, paper_tilemap
  403=>x"17B0",	-- 0001011110110000  
  404=>x"0AEB",	-- 0000101011101011  sub	r3, r5, r3
  405=>x"6E20",	-- 0110111000100000  shr	r0, r4, 7
  406=>x"6219",	-- 0110001000011001  shr	r1, r3, 1
  407=>x"4409",	-- 0100010000001001  shl	r1, r1, 2
  408=>x"C0DA",	-- 1100000011011010  li	r2, 27
  409=>x"0889",	-- 0000100010001001  add	r1, r1, r2
  410=>x"FFF2",	-- 1111111111110010  liw	r2, paper_pos + 1
  411=>x"179E",	-- 0001011110011110  
  412=>x"D012",	-- 1101000000010010  lw	r2, r2
  413=>x"6412",	-- 0110010000010010  shr	r2, r2, 2
  414=>x"C03B",	-- 1100000000111011  li	r3, 7
  415=>x"20D2",	-- 0010000011010010  and	r2, r2, r3
  416=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  417=>x"4E24",	-- 0100111000100100  shl	r4, r4, 7
  418=>x"6E24",	-- 0110111000100100  shr	r4, r4, 7
  419=>x"C00B",	-- 1100000000001011  li	r3, 1
  420=>x"FB06",	-- 1111101100000110  bailne	r0, r6, put_tile
  421=>x"0237",	-- 0000001000110111  
  422=>x"C013",	-- 1100000000010011  li	r3, 2
  423=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_tile
  424=>x"0237",	-- 0000001000110111  
  425=>x"0624",	-- 0000011000100100  dec	r4, r4
  426=>x"BF64",	-- 1011111101100100  brine	r4, PaperGameSegmentLoop
  427=>x"C003",	-- 1100000000000011  li	r3, 0
  428=>x"C144",	-- 1100000101000100  li	r4, 40
  429=>x"0B04",	-- 0000101100000100  sub	r4, r0, r4
  430=>x"FB66",	-- 1111101101100110  baillt	r4, r6, put_tile
  431=>x"0237",	-- 0000001000110111  
  432=>x"D03D",	-- 1101000000111101  lw	r5, r7
  433=>x"043F",	-- 0000010000111111  inc	r7, r7
  434=>x"FFF4",	-- 1111111111110100  liw r4, paper_tilemap + 125
  435=>x"182D",	-- 0001100000101101  
  436=>x"0B2C",	-- 0000101100101100  sub	r4, r5, r4
  437=>x"B625",	-- 1011011000100101  brilt	r4, PaperGameTileLoop
  438=>x"FFF3",	-- 1111111111110011  liw	r3, paper_speed
  439=>x"17A0",	-- 0001011110100000  
  440=>x"D01B",	-- 1101000000011011  lw	r3, r3
  441=>x"CFC4",	-- 1100111111000100  li	r4, 0x1F8
  442=>x"211C",	-- 0010000100011100  and	r4, r3, r4
  443=>x"0924",	-- 0000100100100100  add	r4, r4, r4
  444=>x"0924",	-- 0000100100100100  add	r4, r4, r4
  445=>x"FFF3",	-- 1111111111110011  liw	r3, paper_pos
  446=>x"179D",	-- 0001011110011101  
  447=>x"D018",	-- 1101000000011000  lw	r0, r3
  448=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  449=>x"FFF2",	-- 1111111111110010  liw	r2, paper_sprites
  450=>x"1720",	-- 0001011100100000  
  451=>x"0912",	-- 0000100100010010  add	r2, r2, r4
  452=>x"C161",	-- 1100000101100001  li	r1, 44
  453=>x"C083",	-- 1100000010000011  li	r3, 16
  454=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_16_masked
  455=>x"02FF",	-- 0000001011111111  
  456=>x"92EC",	-- 1001001011101100  brine	r5, PaperGameFail
  458=>x"C028",	-- 1100000000101000  li	r0, 5
  459=>x"C001",	-- 1100000000000001  li	r1, 0
  460=>x"8043",	-- 1000000001000011  bri	-, $+1
  461=>x"8043",	-- 1000000001000011  bri	-, $+1
  462=>x"0609",	-- 0000011000001001  dec	r1, r1
  463=>x"BF4C",	-- 1011111101001100  brine	r1, $-3
  464=>x"0600",	-- 0000011000000000  dec	r0, r0
  465=>x"BE84",	-- 1011111010000100  brine	r0, $-6
  466=>x"FFF2",	-- 1111111111110010  liw	r2, paper_pos
  467=>x"179D",	-- 0001011110011101  
  468=>x"FFF3",	-- 1111111111110011  liw	r3, paper_speed
  469=>x"17A0",	-- 0001011110100000  
  470=>x"D010",	-- 1101000000010000  lw	r0, r2
  471=>x"D019",	-- 1101000000011001  lw	r1, r3
  472=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  473=>x"8E85",	-- 1000111010000101  brilt	r0, PaperGameFail
  474=>x"FFF4",	-- 1111111111110100  liw	r4, 300*8
  475=>x"0960",	-- 0000100101100000  
  476=>x"0B04",	-- 0000101100000100  sub	r4, r0, r4
  477=>x"8DA1",	-- 1000110110100001  brige	r4, PaperGameFail
  478=>x"D210",	-- 1101001000010000  sw	r0, r2
  479=>x"0412",	-- 0000010000010010  inc	r2, r2
  480=>x"041B",	-- 0000010000011011  inc	r3, r3
  481=>x"D010",	-- 1101000000010000  lw	r0, r2
  482=>x"D019",	-- 1101000000011001  lw	r1, r3
  483=>x"C1FC",	-- 1100000111111100  li	r4, 0x3F
  484=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  485=>x"2101",	-- 0010000100000001  and	r1, r0, r4
  486=>x"2624",	-- 0010011000100100  not	r4, r4
  487=>x"2100",	-- 0010000100000000  and	r0, r0, r4
  488=>x"D211",	-- 1101001000010001  sw	r1, r2
  489=>x"83C0",	-- 1000001111000000  brieq	r0, PaperGameSkipScroll
  490=>x"FFF0",	-- 1111111111110000  liw	r0, paper_tilemap
  491=>x"17B0",	-- 0001011110110000  
  492=>x"C021",	-- 1100000000100001  li	r1, 4
  493=>x"0841",	-- 0000100001000001  add	r1, r0, r1
  494=>x"C302",	-- 1100001100000010  li	r2, 24*4
  495=>x"D00B",	-- 1101000000001011  lw	r3, r1
  496=>x"D203",	-- 1101001000000011  sw	r3, r0
  497=>x"0400",	-- 0000010000000000  inc	r0, r0
  498=>x"0409",	-- 0000010000001001  inc	r1, r1
  499=>x"0612",	-- 0000011000010010  dec	r2, r2
  500=>x"BED4",	-- 1011111011010100  brine	r2, PaperGameScrollLoop
  501=>x"C111",	-- 1100000100010001  li	r1, 34
  502=>x"D201",	-- 1101001000000001  sw	r1, r0
  503=>x"0400",	-- 0000010000000000  inc	r0, r0
  504=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  505=>x"16C0",	-- 0001011011000000  
  506=>x"D01B",	-- 1101000000011011  lw	r3, r3
  507=>x"F818",	-- 1111100000011000  baieq	r3, PaperGameRedrawContent
  508=>x"0182",	-- 0000000110000010  
  509=>x"F7DC",	-- 1111011111011100  bspl	r4, r3, 15
  510=>x"88A4",	-- 1000100010100100  brine	r4, PaperGameQuit
  511=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  512=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveUp
  513=>x"F49C",	-- 1111010010011100  bspl	r4, r3, 2
  514=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveDOWN
  515=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  516=>x"81A0",	-- 1000000110100000  brieq	r4, PaperNoMoveLEFT
  517=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  518=>x"17A0",	-- 0001011110100000  
  519=>x"D010",	-- 1101000000010000  lw	r0, r2
  520=>x"0600",	-- 0000011000000000  dec	r0, r0
  521=>x"D210",	-- 1101001000010000  sw	r0, r2
  522=>x"F4DC",	-- 1111010011011100  bspl	r4, r3, 3
  523=>x"81A0",	-- 1000000110100000  brieq	r4, PaperNoMoveRIGHT
  524=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  525=>x"17A0",	-- 0001011110100000  
  526=>x"D010",	-- 1101000000010000  lw	r0, r2
  527=>x"0400",	-- 0000010000000000  inc	r0, r0
  528=>x"D210",	-- 1101001000010000  sw	r0, r2
  529=>x"F8C0",	-- 1111100011000000  bai	-, PaperGameRedrawContent
  530=>x"0182",	-- 0000000110000010  
  531=>x"C000",	-- 1100000000000000  li	r0, 0
  532=>x"FFF2",	-- 1111111111110010  liw	r2, 240*20
  533=>x"12C0",	-- 0001001011000000  
  534=>x"D001",	-- 1101000000000001  lw	r1, r0
  535=>x"2609",	-- 0010011000001001  not	r1, r1
  536=>x"D201",	-- 1101001000000001  sw	r1, r0
  537=>x"0400",	-- 0000010000000000  inc	r0, r0
  538=>x"0612",	-- 0000011000010010  dec	r2, r2
  539=>x"BED4",	-- 1011111011010100  brine	r2, $-5
  540=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  541=>x"16C0",	-- 0001011011000000  
  542=>x"D01A",	-- 1101000000011010  lw	r2, r3
  543=>x"BFD0",	-- 1011111111010000  brieq	r2, $-1
  544=>x"FFFF",	-- 1111111111111111  reset
  545=>x"FFF2",	-- 1111111111110010  liw	r2, rand_seed
  546=>x"16C8",	-- 0001011011001000  
  547=>x"D210",	-- 1101001000010000  sw	r0, r2
  548=>x"E383",	-- 1110001110000011  ba	-, r6
  549=>x"FFF2",	-- 1111111111110010  liw	r2, rand_seed
  550=>x"16C8",	-- 0001011011001000  
  551=>x"D013",	-- 1101000000010011  lw	r3, r2
  552=>x"C7EC",	-- 1100011111101100  li	r4, 253
  553=>x"1F19",	-- 0001111100011001  mixll	r1, r3, r4
  554=>x"18E4",	-- 0001100011100100  mixhh	r4, r4, r3
  555=>x"C002",	-- 1100000000000010  li	r2, 0
  556=>x"0AC9",	-- 0000101011001001  sub	r1, r1, r3
  557=>x"0EA4",	-- 0000111010100100  sbc	r4, r4, r2
  558=>x"0EC9",	-- 0000111011001001  sbc	r1, r1, r3
  559=>x"0EA4",	-- 0000111010100100  sbc	r4, r4, r2
  560=>x"1B13",	-- 0001101100010011  mixhl	r3, r2, r4
  561=>x"0EC9",	-- 0000111011001001  sbc	r1, r1, r3
  562=>x"0C89",	-- 0000110010001001  adc	r1, r1, r2
  563=>x"FFF2",	-- 1111111111110010  liw	r2, rand_seed
  564=>x"16C8",	-- 0001011011001000  
  565=>x"D211",	-- 1101001000010001  sw	r1, r2
  566=>x"E383",	-- 1110001110000011  ba	-, r6
  567=>x"063F",	-- 0000011000111111  dec	r7, r7
  568=>x"D238",	-- 1101001000111000  sw	r0, r7
  569=>x"063F",	-- 0000011000111111  dec	r7, r7
  570=>x"D239",	-- 1101001000111001  sw	r1, r7
  571=>x"063F",	-- 0000011000111111  dec	r7, r7
  572=>x"D23A",	-- 1101001000111010  sw	r2, r7
  573=>x"063F",	-- 0000011000111111  dec	r7, r7
  574=>x"D23B",	-- 1101001000111011  sw	r3, r7
  575=>x"063F",	-- 0000011000111111  dec	r7, r7
  576=>x"D23C",	-- 1101001000111100  sw	r4, r7
  577=>x"063F",	-- 0000011000111111  dec	r7, r7
  578=>x"D23D",	-- 1101001000111101  sw	r5, r7
  579=>x"063F",	-- 0000011000111111  dec	r7, r7
  580=>x"D23E",	-- 1101001000111110  sw	r6, r7
  581=>x"FFF2",	-- 1111111111110010  liw	r2, paper_tiles
  582=>x"1790",	-- 0001011110010000  
  583=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  584=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  585=>x"C043",	-- 1100000001000011  li	r3, 8
  586=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  587=>x"0330",	-- 0000001100110000  
  588=>x"D03E",	-- 1101000000111110  lw	r6, r7
  589=>x"043F",	-- 0000010000111111  inc	r7, r7
  590=>x"D03D",	-- 1101000000111101  lw	r5, r7
  591=>x"043F",	-- 0000010000111111  inc	r7, r7
  592=>x"D03C",	-- 1101000000111100  lw	r4, r7
  593=>x"043F",	-- 0000010000111111  inc	r7, r7
  594=>x"D03B",	-- 1101000000111011  lw	r3, r7
  595=>x"043F",	-- 0000010000111111  inc	r7, r7
  596=>x"D03A",	-- 1101000000111010  lw	r2, r7
  597=>x"043F",	-- 0000010000111111  inc	r7, r7
  598=>x"D039",	-- 1101000000111001  lw	r1, r7
  599=>x"043F",	-- 0000010000111111  inc	r7, r7
  600=>x"D038",	-- 1101000000111000  lw	r0, r7
  601=>x"043F",	-- 0000010000111111  inc	r7, r7
  602=>x"0400",	-- 0000010000000000  inc	r0, r0
  603=>x"E383",	-- 1110001110000011  ba	-, r6
  604=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  605=>x"C084",	-- 1100000010000100  li	r4, 16
  606=>x"0800",	-- 0000100000000000  add	r0, r0, r0
  607=>x"0C49",	-- 0000110001001001  adc	r1, r1, r1
  608=>x"0A8B",	-- 0000101010001011  sub	r3, r1, r2
  609=>x"80DD",	-- 1000000011011101  brilt	r3, div_16_16.skip
  610=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  611=>x"0400",	-- 0000010000000000  inc	r0, r0
  612=>x"0624",	-- 0000011000100100  dec	r4, r4
  613=>x"BE64",	-- 1011111001100100  brine	r4, div_16_16.loop
  614=>x"E383",	-- 1110001110000011  ba	-, r6
  615=>x"063F",	-- 0000011000111111  dec	r7, r7
  616=>x"D23E",	-- 1101001000111110  sw	r6, r7
  617=>x"D013",	-- 1101000000010011  lw	r3, r2
  618=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  619=>x"84D8",	-- 1000010011011000  brieq	r3, puts.end
  620=>x"063F",	-- 0000011000111111  dec	r7, r7
  621=>x"D23A",	-- 1101001000111010  sw	r2, r7
  622=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  623=>x"0281",	-- 0000001010000001  
  624=>x"D03A",	-- 1101000000111010  lw	r2, r7
  625=>x"043F",	-- 0000010000111111  inc	r7, r7
  626=>x"D013",	-- 1101000000010011  lw	r3, r2
  627=>x"4E1B",	-- 0100111000011011  shl	r3, r3, 7
  628=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  629=>x"8258",	-- 1000001001011000  brieq	r3, puts.end
  630=>x"063F",	-- 0000011000111111  dec	r7, r7
  631=>x"D23A",	-- 1101001000111010  sw	r2, r7
  632=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  633=>x"0281",	-- 0000001010000001  
  634=>x"D03A",	-- 1101000000111010  lw	r2, r7
  635=>x"043F",	-- 0000010000111111  inc	r7, r7
  636=>x"0412",	-- 0000010000010010  inc	r2, r2
  637=>x"BB03",	-- 1011101100000011  bri	-, puts.loop
  638=>x"D03E",	-- 1101000000111110  lw	r6, r7
  639=>x"043F",	-- 0000010000111111  inc	r7, r7
  640=>x"E383",	-- 1110001110000011  ba	-, r6
  641=>x"063F",	-- 0000011000111111  dec	r7, r7
  642=>x"D23E",	-- 1101001000111110  sw	r6, r7
  643=>x"063F",	-- 0000011000111111  dec	r7, r7
  644=>x"D238",	-- 1101001000111000  sw	r0, r7
  645=>x"063F",	-- 0000011000111111  dec	r7, r7
  646=>x"D239",	-- 1101001000111001  sw	r1, r7
  647=>x"FFF2",	-- 1111111111110010  liw	r2, font_map
  648=>x"12C0",	-- 0001001011000000  
  649=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  650=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  651=>x"C043",	-- 1100000001000011  li	r3, 8
  652=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  653=>x"0330",	-- 0000001100110000  
  654=>x"D039",	-- 1101000000111001  lw	r1, r7
  655=>x"043F",	-- 0000010000111111  inc	r7, r7
  656=>x"D038",	-- 1101000000111000  lw	r0, r7
  657=>x"043F",	-- 0000010000111111  inc	r7, r7
  658=>x"0400",	-- 0000010000000000  inc	r0, r0
  659=>x"D03E",	-- 1101000000111110  lw	r6, r7
  660=>x"043F",	-- 0000010000111111  inc	r7, r7
  661=>x"E383",	-- 1110001110000011  ba	-, r6
  662=>x"063F",	-- 0000011000111111  dec	r7, r7
  663=>x"D23E",	-- 1101001000111110  sw	r6, r7
  664=>x"FFF4",	-- 1111111111110100  liw	r4, 10000
  665=>x"2710",	-- 0010011100010000  
  666=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  667=>x"02A9",	-- 0000001010101001  
  668=>x"FFF4",	-- 1111111111110100  liw	r4, 1000
  669=>x"03E8",	-- 0000001111101000  
  670=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  671=>x"02A9",	-- 0000001010101001  
  672=>x"C324",	-- 1100001100100100  li	r4, 100
  673=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  674=>x"02A9",	-- 0000001010101001  
  675=>x"C054",	-- 1100000001010100  li	r4, 10
  676=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  677=>x"02A9",	-- 0000001010101001  
  678=>x"D03E",	-- 1101000000111110  lw	r6, r7
  679=>x"043F",	-- 0000010000111111  inc	r7, r7
  680=>x"C00C",	-- 1100000000001100  li	r4, 1
  681=>x"C17B",	-- 1100000101111011  li	r3, 0x2F
  682=>x"041B",	-- 0000010000011011  inc	r3, r3
  683=>x"0B12",	-- 0000101100010010  sub	r2, r2, r4
  684=>x"BF91",	-- 1011111110010001  brige	r2, printnum.loop
  685=>x"0912",	-- 0000100100010010  add	r2, r2, r4
  686=>x"063F",	-- 0000011000111111  dec	r7, r7
  687=>x"D23E",	-- 1101001000111110  sw	r6, r7
  688=>x"063F",	-- 0000011000111111  dec	r7, r7
  689=>x"D23A",	-- 1101001000111010  sw	r2, r7
  690=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  691=>x"0281",	-- 0000001010000001  
  692=>x"D03A",	-- 1101000000111010  lw	r2, r7
  693=>x"043F",	-- 0000010000111111  inc	r7, r7
  694=>x"D03E",	-- 1101000000111110  lw	r6, r7
  695=>x"043F",	-- 0000010000111111  inc	r7, r7
  696=>x"E383",	-- 1110001110000011  ba	-, r6
  697=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  698=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  699=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  700=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  701=>x"C0A0",	-- 1100000010100000  li	r0, 20
  702=>x"D011",	-- 1101000000010001  lw	r1, r2
  703=>x"D221",	-- 1101001000100001  sw	r1, r4
  704=>x"0412",	-- 0000010000010010  inc	r2, r2
  705=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  706=>x"061B",	-- 0000011000011011  dec	r3, r3
  707=>x"BEDC",	-- 1011111011011100  brine	r3, put_sprite_16_aligned.loop
  708=>x"E383",	-- 1110001110000011  ba	-, r6
  709=>x"C07D",	-- 1100000001111101  li	r5, 15
  710=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  711=>x"6600",	-- 0110011000000000  shr	r0, r0, 3
  712=>x"BC68",	-- 1011110001101000  brieq	r5, put_sprite_16_aligned
  713=>x"062D",	-- 0000011000101101  dec	r5, r5
  714=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  715=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  716=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  717=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  718=>x"063F",	-- 0000011000111111  dec	r7, r7
  719=>x"D23B",	-- 1101001000111011  sw	r3, r7
  720=>x"D011",	-- 1101000000010001  lw	r1, r2
  721=>x"CFF8",	-- 1100111111111000  li	r0, -1
  722=>x"3D40",	-- 0011110101000000  rsr	r0, r0, r5
  723=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  724=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  725=>x"D023",	-- 1101000000100011  lw	r3, r4
  726=>x"2600",	-- 0010011000000000  not	r0, r0
  727=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  728=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  729=>x"D221",	-- 1101001000100001  sw	r1, r4
  730=>x"0424",	-- 0000010000100100  inc	r4, r4
  731=>x"D011",	-- 1101000000010001  lw	r1, r2
  732=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  733=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  734=>x"D023",	-- 1101000000100011  lw	r3, r4
  735=>x"2600",	-- 0010011000000000  not	r0, r0
  736=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  737=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  738=>x"D221",	-- 1101001000100001  sw	r1, r4
  739=>x"0412",	-- 0000010000010010  inc	r2, r2
  740=>x"C098",	-- 1100000010011000  li	r0, 19
  741=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  742=>x"D03B",	-- 1101000000111011  lw	r3, r7
  743=>x"043F",	-- 0000010000111111  inc	r7, r7
  744=>x"061B",	-- 0000011000011011  dec	r3, r3
  745=>x"B95C",	-- 1011100101011100  brine	r3, put_sprite_16.loop
  746=>x"E383",	-- 1110001110000011  ba	-, r6
  747=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  748=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  749=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  750=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  751=>x"C005",	-- 1100000000000101  li	r5, 0
  752=>x"D020",	-- 1101000000100000  lw	r0, r4
  753=>x"D011",	-- 1101000000010001  lw	r1, r2
  754=>x"0412",	-- 0000010000010010  inc	r2, r2
  755=>x"2040",	-- 0010000001000000  and	r0, r0, r1
  756=>x"D011",	-- 1101000000010001  lw	r1, r2
  757=>x"0412",	-- 0000010000010010  inc	r2, r2
  758=>x"2240",	-- 0010001001000000  or	r0, r0, r1
  759=>x"E420",	-- 1110010000100000  exw	r0, r4
  760=>x"2040",	-- 0010000001000000  and	r0, r0, r1
  761=>x"222D",	-- 0010001000101101  or	r5, r5, r0
  762=>x"C0A0",	-- 1100000010100000  li	r0, 20
  763=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  764=>x"061B",	-- 0000011000011011  dec	r3, r3
  765=>x"B05C",	-- 1011000001011100  brine	r3, put_sprite_16_aligned.loop
  766=>x"E383",	-- 1110001110000011  ba	-, r6
  767=>x"C07D",	-- 1100000001111101  li	r5, 15
  768=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  769=>x"6600",	-- 0110011000000000  shr	r0, r0, 3
  770=>x"BA68",	-- 1011101001101000  brieq	r5, put_sprite_16_masked_aligned
  771=>x"062D",	-- 0000011000101101  dec	r5, r5
  772=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  773=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  774=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  775=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  776=>x"063F",	-- 0000011000111111  dec	r7, r7
  777=>x"D23E",	-- 1101001000111110  sw	r6, r7
  778=>x"102E",	-- 0001000000101110  mova	r6, r5
  779=>x"C005",	-- 1100000000000101  li	r5, 0
  780=>x"063F",	-- 0000011000111111  dec	r7, r7
  781=>x"D23B",	-- 1101001000111011  sw	r3, r7
  782=>x"D010",	-- 1101000000010000  lw	r0, r2
  783=>x"0412",	-- 0000010000010010  inc	r2, r2
  784=>x"3D80",	-- 0011110110000000  rsr	r0, r0, r6
  785=>x"D011",	-- 1101000000010001  lw	r1, r2
  786=>x"3989",	-- 0011100110001001  rrr	r1, r1, r6
  787=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  788=>x"D023",	-- 1101000000100011  lw	r3, r4
  789=>x"2600",	-- 0010011000000000  not	r0, r0
  790=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  791=>x"225B",	-- 0010001001011011  or	r3, r3, r1
  792=>x"E423",	-- 1110010000100011  exw	r3, r4
  793=>x"205B",	-- 0010000001011011  and	r3, r3, r1
  794=>x"22ED",	-- 0010001011101101  or	r5, r5, r3
  795=>x"0424",	-- 0000010000100100  inc	r4, r4
  796=>x"D011",	-- 1101000000010001  lw	r1, r2
  797=>x"3989",	-- 0011100110001001  rrr	r1, r1, r6
  798=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  799=>x"D023",	-- 1101000000100011  lw	r3, r4
  800=>x"2600",	-- 0010011000000000  not	r0, r0
  801=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  802=>x"225B",	-- 0010001001011011  or	r3, r3, r1
  803=>x"E423",	-- 1110010000100011  exw	r3, r4
  804=>x"205B",	-- 0010000001011011  and	r3, r3, r1
  805=>x"22ED",	-- 0010001011101101  or	r5, r5, r3
  806=>x"0412",	-- 0000010000010010  inc	r2, r2
  807=>x"C098",	-- 1100000010011000  li	r0, 19
  808=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  809=>x"D03B",	-- 1101000000111011  lw	r3, r7
  810=>x"043F",	-- 0000010000111111  inc	r7, r7
  811=>x"061B",	-- 0000011000011011  dec	r3, r3
  812=>x"B81C",	-- 1011100000011100  brine	r3, put_sprite_16_masked.loop
  813=>x"D03E",	-- 1101000000111110  lw	r6, r7
  814=>x"043F",	-- 0000010000111111  inc	r7, r7
  815=>x"E383",	-- 1110001110000011  ba	-, r6
  816=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  817=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  818=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  819=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  820=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  821=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  822=>x"C0A5",	-- 1100000010100101  li	r5, 20
  823=>x"8404",	-- 1000010000000100  brine	r0, put_sprite_8_aligned.loop1
  824=>x"D010",	-- 1101000000010000  lw	r0, r2
  825=>x"D021",	-- 1101000000100001  lw	r1, r4
  826=>x"1A41",	-- 0001101001000001  mixhl	r1, r0, r1
  827=>x"D221",	-- 1101001000100001  sw	r1, r4
  828=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  829=>x"061B",	-- 0000011000011011  dec	r3, r3
  830=>x"E398",	-- 1110001110011000  baeq	r3, r6
  831=>x"D021",	-- 1101000000100001  lw	r1, r4
  832=>x"1E41",	-- 0001111001000001  mixll	r1, r0, r1
  833=>x"D221",	-- 1101001000100001  sw	r1, r4
  834=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  835=>x"0412",	-- 0000010000010010  inc	r2, r2
  836=>x"061B",	-- 0000011000011011  dec	r3, r3
  837=>x"E398",	-- 1110001110011000  baeq	r3, r6
  838=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop0
  839=>x"D010",	-- 1101000000010000  lw	r0, r2
  840=>x"D021",	-- 1101000000100001  lw	r1, r4
  841=>x"1809",	-- 0001100000001001  mixhh	r1, r1, r0
  842=>x"D221",	-- 1101001000100001  sw	r1, r4
  843=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  844=>x"061B",	-- 0000011000011011  dec	r3, r3
  845=>x"E398",	-- 1110001110011000  baeq	r3, r6
  846=>x"D021",	-- 1101000000100001  lw	r1, r4
  847=>x"1A09",	-- 0001101000001001  mixhl	r1, r1, r0
  848=>x"D221",	-- 1101001000100001  sw	r1, r4
  849=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  850=>x"0412",	-- 0000010000010010  inc	r2, r2
  851=>x"061B",	-- 0000011000011011  dec	r3, r3
  852=>x"E398",	-- 1110001110011000  baeq	r3, r6
  853=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop1
  854=>x"C03D",	-- 1100000000111101  li	r5, 7
  855=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  856=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  857=>x"B5E8",	-- 1011010111101000  brieq	r5, put_sprite_8_aligned
  858=>x"062D",	-- 0000011000101101  dec	r5, r5
  859=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  860=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  861=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  862=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  863=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  864=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  865=>x"8A04",	-- 1000101000000100  brine	r0, put_sprite_8.loop1
  866=>x"D010",	-- 1101000000010000  lw	r0, r2
  867=>x"063F",	-- 0000011000111111  dec	r7, r7
  868=>x"D23A",	-- 1101001000111010  sw	r2, r7
  869=>x"C802",	-- 1100100000000010  li	r2, 0x100
  870=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  871=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  872=>x"D021",	-- 1101000000100001  lw	r1, r4
  873=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  874=>x"2612",	-- 0010011000010010  not	r2, r2
  875=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  876=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  877=>x"D221",	-- 1101001000100001  sw	r1, r4
  878=>x"C0A1",	-- 1100000010100001  li	r1, 20
  879=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  880=>x"D03A",	-- 1101000000111010  lw	r2, r7
  881=>x"043F",	-- 0000010000111111  inc	r7, r7
  882=>x"061B",	-- 0000011000011011  dec	r3, r3
  883=>x"E398",	-- 1110001110011000  baeq	r3, r6
  884=>x"D010",	-- 1101000000010000  lw	r0, r2
  885=>x"063F",	-- 0000011000111111  dec	r7, r7
  886=>x"D23A",	-- 1101001000111010  sw	r2, r7
  887=>x"1E00",	-- 0001111000000000  mixll	r0, r0, r0
  888=>x"C802",	-- 1100100000000010  li	r2, 0x100
  889=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  890=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  891=>x"D021",	-- 1101000000100001  lw	r1, r4
  892=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  893=>x"2612",	-- 0010011000010010  not	r2, r2
  894=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  895=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  896=>x"D221",	-- 1101001000100001  sw	r1, r4
  897=>x"C0A1",	-- 1100000010100001  li	r1, 20
  898=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  899=>x"D03A",	-- 1101000000111010  lw	r2, r7
  900=>x"043F",	-- 0000010000111111  inc	r7, r7
  901=>x"0412",	-- 0000010000010010  inc	r2, r2
  902=>x"061B",	-- 0000011000011011  dec	r3, r3
  903=>x"E398",	-- 1110001110011000  baeq	r3, r6
  904=>x"B683",	-- 1011011010000011  bri	-, put_sprite_8.loop0
  905=>x"D010",	-- 1101000000010000  lw	r0, r2
  906=>x"063F",	-- 0000011000111111  dec	r7, r7
  907=>x"D23A",	-- 1101001000111010  sw	r2, r7
  908=>x"063F",	-- 0000011000111111  dec	r7, r7
  909=>x"D23B",	-- 1101001000111011  sw	r3, r7
  910=>x"C802",	-- 1100100000000010  li	r2, 0x100
  911=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  912=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  913=>x"2080",	-- 0010000010000000  and	r0, r0, r2
  914=>x"D021",	-- 1101000000100001  lw	r1, r4
  915=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
  916=>x"261B",	-- 0010011000011011  not	r3, r3
  917=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  918=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
  919=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  920=>x"D221",	-- 1101001000100001  sw	r1, r4
  921=>x"0424",	-- 0000010000100100  inc	r4, r4
  922=>x"D021",	-- 1101000000100001  lw	r1, r4
  923=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  924=>x"261B",	-- 0010011000011011  not	r3, r3
  925=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  926=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
  927=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  928=>x"D221",	-- 1101001000100001  sw	r1, r4
  929=>x"C099",	-- 1100000010011001  li	r1, 19
  930=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  931=>x"D03B",	-- 1101000000111011  lw	r3, r7
  932=>x"043F",	-- 0000010000111111  inc	r7, r7
  933=>x"D03A",	-- 1101000000111010  lw	r2, r7
  934=>x"043F",	-- 0000010000111111  inc	r7, r7
  935=>x"061B",	-- 0000011000011011  dec	r3, r3
  936=>x"E398",	-- 1110001110011000  baeq	r3, r6
  937=>x"D010",	-- 1101000000010000  lw	r0, r2
  938=>x"4E00",	-- 0100111000000000  shl	r0, r0, 7
  939=>x"063F",	-- 0000011000111111  dec	r7, r7
  940=>x"D23A",	-- 1101001000111010  sw	r2, r7
  941=>x"063F",	-- 0000011000111111  dec	r7, r7
  942=>x"D23B",	-- 1101001000111011  sw	r3, r7
  943=>x"C802",	-- 1100100000000010  li	r2, 0x100
  944=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  945=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  946=>x"2080",	-- 0010000010000000  and	r0, r0, r2
  947=>x"D021",	-- 1101000000100001  lw	r1, r4
  948=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
  949=>x"261B",	-- 0010011000011011  not	r3, r3
  950=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  951=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
  952=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  953=>x"D221",	-- 1101001000100001  sw	r1, r4
  954=>x"0424",	-- 0000010000100100  inc	r4, r4
  955=>x"D021",	-- 1101000000100001  lw	r1, r4
  956=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  957=>x"261B",	-- 0010011000011011  not	r3, r3
  958=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  959=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
  960=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  961=>x"D221",	-- 1101001000100001  sw	r1, r4
  962=>x"C099",	-- 1100000010011001  li	r1, 19
  963=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  964=>x"D03B",	-- 1101000000111011  lw	r3, r7
  965=>x"043F",	-- 0000010000111111  inc	r7, r7
  966=>x"D03A",	-- 1101000000111010  lw	r2, r7
  967=>x"043F",	-- 0000010000111111  inc	r7, r7
  968=>x"0412",	-- 0000010000010010  inc	r2, r2
  969=>x"061B",	-- 0000011000011011  dec	r3, r3
  970=>x"E398",	-- 1110001110011000  baeq	r3, r6
  971=>x"AF83",	-- 1010111110000011  bri	-, put_sprite_8.loop1
    others => x"0000"
    );
begin
  process(CLK)
  begin
    if (CLK'event AND CLK='1') then
      D <= m(to_integer(unsigned(AD)));
    end if;
  end process;
end Behavioral;
