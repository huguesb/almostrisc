----------------------------------------------------------------------------------
--
-- File retrieved, on 07/02/2010, from :
-- http://sebastien-viardot.imag.fr/Enseignements/Archi1A2s/sources/ROMPROG.vhd
--
-- Slightly altered to get rid of vendor-specific packages and adjust formatting
-- Now auto-filled by asrom script
--
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROMPROG is
  Port ( AD : in  STD_LOGIC_VECTOR (12 downto 0);
         D : out  STD_LOGIC_VECTOR (15 downto 0);
         CLK : in STD_LOGIC);
end ROMPROG;

architecture Behavioral of ROMPROG is
  constant low_address: natural := 0;
  constant high_address: natural := 8192;
  subtype octet is std_logic_vector( 15 downto 0 );
  type zone_memoire is
    array (natural range low_address to high_address-1) of octet;
  constant m: zone_memoire:= (
    0=>x"FFF7",	-- 1111111111110111  liw	r7, IRQ_mask
    1=>x"2000",	-- 0010000000000000  
    2=>x"F8C0",	-- 1111100011000000  bai	-, os_init
    3=>x"0100",	-- 0000000100000000  
   16=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_ack
   17=>x"2002",	-- 0010000000000010  
   18=>x"D001",	-- 1101000000000001  lw	r1, r0
   19=>x"F54A",	-- 1111010101001010  bspl	r2, r1, 5
   20=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_error
   21=>x"0050",	-- 0000000001010000  
   22=>x"F4CA",	-- 1111010011001010  bspl	r2, r1, 3
   23=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_kbd
   24=>x"0060",	-- 0000000001100000  
   25=>x"F40A",	-- 1111010000001010  bspl	r2, r1, 0
   26=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_tmr
   27=>x"0040",	-- 0000000001000000  
   28=>x"D201",	-- 1101001000000001  sw	r1, r0
   29=>x"FFFE",	-- 1111111111111110  reti
   64=>x"263F",	-- 0010011000111111  not r7, r7
   65=>x"D7C0",	-- 1101011111000000  out	r7
   66=>x"E383",	-- 1110001110000011  ba	-, r6
   80=>x"25FF",	-- 0010010111111111  xor	r7, r7, r7
   81=>x"D7C0",	-- 1101011111000000  out	r7
   82=>x"E383",	-- 1110001110000011  ba	-, r6
   96=>x"FFF2",	-- 1111111111110010  liw	r2, PS2_rx
   97=>x"2004",	-- 0010000000000100  
   98=>x"D012",	-- 1101000000010010  lw	r2, r2
   99=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map + 8
  100=>x"1808",	-- 0001100000001000  
  101=>x"D01B",	-- 1101000000011011  lw	r3, r3
  102=>x"1EBF",	-- 0001111010111111  mixll	r7, r7, r2
  103=>x"C784",	-- 1100011110000100  li	r4, 0xF0
  104=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  105=>x"8B20",	-- 1000101100100000  brieq	r4, int_kbd.release
  106=>x"C704",	-- 1100011100000100  li	r4, 0xE0
  107=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  108=>x"88E0",	-- 1000100011100000  brieq	r4, int_kbd.extended
  109=>x"FFF5",	-- 1111111111110101  liw	r5, paper_keys - 1
  110=>x"16BF",	-- 0001011010111111  
  111=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  112=>x"80E0",	-- 1000000011100000  brieq	r4, $+3
  113=>x"FFF5",	-- 1111111111110101  liw	r5, paper_keys + 11 - 1
  114=>x"16CA",	-- 0001011011001010  
  115=>x"042D",	-- 0000010000101101  inc	r5, r5
  116=>x"D02C",	-- 1101000000101100  lw	r4, r5
  117=>x"8560",	-- 1000010101100000  brieq	r4, scan_code_mismatch
  118=>x"6E24",	-- 0110111000100100  shr	r4, r4, 7
  119=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  120=>x"BEE4",	-- 1011111011100100  brine	r4, scan_code_loop
  121=>x"D02A",	-- 1101000000101010  lw	r2, r5
  122=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  123=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  124=>x"741B",	-- 0111010000011011  shr	r3, r3, 10
  125=>x"C00D",	-- 1100000000001101  li	r5, 1
  126=>x"0612",	-- 0000011000010010  dec	r2, r2
  127=>x"3AAA",	-- 0011101010101010  rrl	r2, r5, r2
  128=>x"FFF5",	-- 1111111111110101  liw	r5, key_press_map
  129=>x"1800",	-- 0001100000000000  
  130=>x"08ED",	-- 0000100011101101  add	r5, r5, r3
  131=>x"D02B",	-- 1101000000101011  lw	r3, r5
  132=>x"80E4",	-- 1000000011100100  brine	r4, scan_code_release
  133=>x"229B",	-- 0010001010011011  or	r3, r3, r2
  134=>x"80C3",	-- 1000000011000011  bri	-, scan_code_notify
  135=>x"2612",	-- 0010011000010010  not	r2, r2
  136=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  137=>x"D22B",	-- 1101001000101011  sw	r3, r5
  138=>x"C003",	-- 1100000000000011  li	r3, 0
  139=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  140=>x"1808",	-- 0001100000001000  
  141=>x"D223",	-- 1101001000100011  sw	r3, r4
  142=>x"E383",	-- 1110001110000011  ba	-, r6
  143=>x"C014",	-- 1100000000010100  li	r4, 2
  144=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  145=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  146=>x"1808",	-- 0001100000001000  
  147=>x"D223",	-- 1101001000100011  sw	r3, r4
  148=>x"E383",	-- 1110001110000011  ba	-, r6
  149=>x"C00C",	-- 1100000000001100  li	r4, 1
  150=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  151=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  152=>x"1808",	-- 0001100000001000  
  153=>x"D223",	-- 1101001000100011  sw	r3, r4
  154=>x"E383",	-- 1110001110000011  ba	-, r6
  256=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_mask
  257=>x"2000",	-- 0010000000000000  
  258=>x"C0C9",	-- 1100000011001001  li	r1, 0x19
  259=>x"D201",	-- 1101001000000001  sw	r1, r0
  260=>x"0400",	-- 0000010000000000  inc	r0, r0
  261=>x"CFF9",	-- 1100111111111001  li	r1, -1
  262=>x"D201",	-- 1101001000000001  sw	r1, r0
  263=>x"C03A",	-- 1100000000111010  li	r2, 7
  264=>x"0880",	-- 0000100010000000  add	r0, r0, r2
  265=>x"C0EA",	-- 1100000011101010  li	r2, 0x1D
  266=>x"D202",	-- 1101001000000010  sw	r2, r0
  267=>x"0400",	-- 0000010000000000  inc	r0, r0
  268=>x"C07A",	-- 1100000001111010  li	r2, 15
  269=>x"D202",	-- 1101001000000010  sw	r2, r0
  270=>x"FFF0",	-- 1111111111110000  liw	r0, key_press_map
  271=>x"1800",	-- 0001100000000000  
  272=>x"C001",	-- 1100000000000001  li	r1, 0
  273=>x"C042",	-- 1100000001000010  li	r2, 8
  274=>x"D201",	-- 1101001000000001  sw	r1, r0
  275=>x"0400",	-- 0000010000000000  inc	r0, r0
  276=>x"0612",	-- 0000011000010010  dec	r2, r2
  277=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  278=>x"C0F3",	-- 1100000011110011  li	r3, 30
  279=>x"CFFA",	-- 1100111111111010  li	r2, -1
  280=>x"D21A",	-- 1101001000011010  sw	r2, r3
  281=>x"8083",	-- 1000000010000011  bri	-, PaperGameStart
  282=>x"8003",	-- 1000000000000011  bri	-, PaperMenuLoop
  283=>x"FFF0",	-- 1111111111110000  liw	r0, paper_dir
  284=>x"173C",	-- 0001011100111100  
  285=>x"C001",	-- 1100000000000001  li	r1, 0
  286=>x"D201",	-- 1101001000000001  sw	r1, r0
  287=>x"0400",	-- 0000010000000000  inc	r0, r0
  288=>x"C4C1",	-- 1100010011000001  li	r1, 152
  289=>x"D201",	-- 1101001000000001  sw	r1, r0
  290=>x"0400",	-- 0000010000000000  inc	r0, r0
  291=>x"C001",	-- 1100000000000001  li	r1, 0
  292=>x"D201",	-- 1101001000000001  sw	r1, r0
  293=>x"0400",	-- 0000010000000000  inc	r0, r0
  294=>x"C401",	-- 1100010000000001  li	r1, 128
  295=>x"D201",	-- 1101001000000001  sw	r1, r0
  296=>x"0400",	-- 0000010000000000  inc	r0, r0
  297=>x"C001",	-- 1100000000000001  li	r1, 0
  298=>x"D201",	-- 1101001000000001  sw	r1, r0
  299=>x"0400",	-- 0000010000000000  inc	r0, r0
  300=>x"C0A1",	-- 1100000010100001  li	r1, 20
  301=>x"D201",	-- 1101001000000001  sw	r1, r0
  302=>x"0400",	-- 0000010000000000  inc	r0, r0
  303=>x"C029",	-- 1100000000101001  li	r1, 5
  304=>x"D201",	-- 1101001000000001  sw	r1, r0
  305=>x"0400",	-- 0000010000000000  inc	r0, r0
  306=>x"C000",	-- 1100000000000000  li	r0, 0
  307=>x"CFF9",	-- 1100111111111001  li	r1, -1
  308=>x"C0A2",	-- 1100000010100010  li	r2, 20
  309=>x"D201",	-- 1101001000000001  sw	r1, r0
  310=>x"0400",	-- 0000010000000000  inc	r0, r0
  311=>x"0612",	-- 0000011000010010  dec	r2, r2
  312=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  313=>x"C001",	-- 1100000000000001  li	r1, 0
  314=>x"FFF2",	-- 1111111111110010  liw	r2, 18*20
  315=>x"0168",	-- 0000000101101000  
  316=>x"D201",	-- 1101001000000001  sw	r1, r0
  317=>x"0400",	-- 0000010000000000  inc	r0, r0
  318=>x"0612",	-- 0000011000010010  dec	r2, r2
  319=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  320=>x"CFF9",	-- 1100111111111001  li	r1, -1
  321=>x"C0A2",	-- 1100000010100010  li	r2, 20
  322=>x"D201",	-- 1101001000000001  sw	r1, r0
  323=>x"0400",	-- 0000010000000000  inc	r0, r0
  324=>x"0612",	-- 0000011000010010  dec	r2, r2
  325=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  326=>x"C020",	-- 1100000000100000  li	r0, 4
  327=>x"C029",	-- 1100000000101001  li	r1, 5
  328=>x"FFF2",	-- 1111111111110010  liw	r2, paper_title
  329=>x"1744",	-- 0001011101000100  
  330=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  331=>x"0236",	-- 0000001000110110  
  332=>x"C778",	-- 1100011101111000  li	r0, 239
  333=>x"C009",	-- 1100000000001001  li	r1, 1
  334=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud
  335=>x"1720",	-- 0001011100100000  
  336=>x"C043",	-- 1100000001000011  li	r3, 8
  337=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  338=>x"02E0",	-- 0000001011100000  
  339=>x"C0F8",	-- 1100000011111000  li	r0, 31
  340=>x"C009",	-- 1100000000001001  li	r1, 1
  341=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed + 1
  342=>x"173E",	-- 0001011100111110  
  343=>x"D012",	-- 1101000000010010  lw	r2, r2
  344=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum
  345=>x"0265",	-- 0000001001100101  
  346=>x"C120",	-- 1100000100100000  li	r0, 36
  347=>x"C009",	-- 1100000000001001  li	r1, 1
  348=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  349=>x"174A",	-- 0001011101001010  
  350=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  351=>x"0236",	-- 0000001000110110  
  352=>x"C778",	-- 1100011101111000  li	r0, 239
  353=>x"C051",	-- 1100000001010001  li	r1, 10
  354=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud + 4
  355=>x"1724",	-- 0001011100100100  
  356=>x"C043",	-- 1100000001000011  li	r3, 8
  357=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  358=>x"02E0",	-- 0000001011100000  
  359=>x"C0F8",	-- 1100000011111000  li	r0, 31
  360=>x"C051",	-- 1100000001010001  li	r1, 10
  361=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed + 2
  362=>x"173F",	-- 0001011100111111  
  363=>x"D012",	-- 1101000000010010  lw	r2, r2
  364=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum
  365=>x"0265",	-- 0000001001100101  
  366=>x"C120",	-- 1100000100100000  li	r0, 36
  367=>x"C051",	-- 1100000001010001  li	r1, 10
  368=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  369=>x"174A",	-- 0001011101001010  
  370=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  371=>x"0236",	-- 0000001000110110  
  372=>x"FFF0",	-- 1111111111110000  liw	r0, 20*20
  373=>x"0190",	-- 0000000110010000  
  374=>x"C001",	-- 1100000000000001  li	r1, 0
  375=>x"FFF2",	-- 1111111111110010  liw	r2, 220*20
  376=>x"1130",	-- 0001000100110000  
  377=>x"D201",	-- 1101001000000001  sw	r1, r0
  378=>x"0400",	-- 0000010000000000  inc	r0, r0
  379=>x"0612",	-- 0000011000010010  dec	r2, r2
  380=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  381=>x"FFF5",	-- 1111111111110101  liw	r5, paper_tilemap
  382=>x"1780",	-- 0001011110000000  
  383=>x"D02C",	-- 1101000000101100  lw	r4, r5
  384=>x"042D",	-- 0000010000101101  inc	r5, r5
  385=>x"8720",	-- 1000011100100000  brieq	r4, PaperGameTileSkip
  386=>x"063F",	-- 0000011000111111  dec	r7, r7
  387=>x"D23D",	-- 1101001000111101  sw	r5, r7
  388=>x"FFF3",	-- 1111111111110011  liw	r3, paper_tilemap
  389=>x"1780",	-- 0001011110000000  
  390=>x"0AEB",	-- 0000101011101011  sub	r3, r5, r3
  391=>x"6E20",	-- 0110111000100000  shr	r0, r4, 7
  392=>x"6219",	-- 0110001000011001  shr	r1, r3, 1
  393=>x"4409",	-- 0100010000001001  shl	r1, r1, 2
  394=>x"FFF2",	-- 1111111111110010  liw	r2, paper_pos + 1
  395=>x"1741",	-- 0001011101000001  
  396=>x"D012",	-- 1101000000010010  lw	r2, r2
  397=>x"6412",	-- 0110010000010010  shr	r2, r2, 2
  398=>x"C03B",	-- 1100000000111011  li	r3, 7
  399=>x"20D2",	-- 0010000011010010  and	r2, r2, r3
  400=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  401=>x"4E24",	-- 0100111000100100  shl	r4, r4, 7
  402=>x"6E24",	-- 0110111000100100  shr	r4, r4, 7
  403=>x"C00B",	-- 1100000000001011  li	r3, 1
  404=>x"FB06",	-- 1111101100000110  bailne	r0, r6, put_tile
  405=>x"01E2",	-- 0000000111100010  
  406=>x"C013",	-- 1100000000010011  li	r3, 2
  407=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_tile
  408=>x"01E2",	-- 0000000111100010  
  409=>x"0624",	-- 0000011000100100  dec	r4, r4
  410=>x"BF64",	-- 1011111101100100  brine	r4, PaperGameSegmentLoop
  411=>x"D03D",	-- 1101000000111101  lw	r5, r7
  412=>x"043F",	-- 0000010000111111  inc	r7, r7
  413=>x"FFF4",	-- 1111111111110100  liw r4, paper_tilemap + 125
  414=>x"17FD",	-- 0001011111111101  
  415=>x"0B2C",	-- 0000101100101100  sub	r4, r5, r4
  416=>x"B7E5",	-- 1011011111100101  brilt	r4, PaperGameTileLoop
  417=>x"FFF3",	-- 1111111111110011  liw	r3, paper_speed
  418=>x"173D",	-- 0001011100111101  
  419=>x"D01C",	-- 1101000000011100  lw	r4, r3
  420=>x"6424",	-- 0110010000100100  shr	r4, r4, 2
  421=>x"041B",	-- 0000010000011011  inc	r3, r3
  422=>x"D018",	-- 1101000000011000  lw	r0, r3
  423=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  424=>x"FFF2",	-- 1111111111110010  liw	r2, paper_sprites
  425=>x"16F0",	-- 0001011011110000  
  426=>x"4624",	-- 0100011000100100  shl	r4, r4, 3
  427=>x"0912",	-- 0000100100010010  add	r2, r2, r4
  428=>x"C161",	-- 1100000101100001  li	r1, 44
  429=>x"C083",	-- 1100000010000011  li	r3, 16
  430=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_16
  431=>x"0294",	-- 0000001010010100  
  432=>x"C01A",	-- 1100000000011010  li	r2, 3
  433=>x"C003",	-- 1100000000000011  li	r3, 0
  434=>x"061B",	-- 0000011000011011  dec	r3, r3
  435=>x"BFDC",	-- 1011111111011100  brine	r3, $-1
  436=>x"0612",	-- 0000011000010010  dec	r2, r2
  437=>x"BF14",	-- 1011111100010100  brine	r2, $-4
  438=>x"FFF2",	-- 1111111111110010  liw	r2, paper_pos
  439=>x"1740",	-- 0001011101000000  
  440=>x"FFF3",	-- 1111111111110011  liw	r3, paper_speed
  441=>x"173D",	-- 0001011100111101  
  442=>x"D010",	-- 1101000000010000  lw	r0, r2
  443=>x"D019",	-- 1101000000011001  lw	r1, r3
  444=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  445=>x"8905",	-- 1000100100000101  brilt	r0, PaperGameQuit
  446=>x"C964",	-- 1100100101100100  li	r4, 300
  447=>x"0B04",	-- 0000101100000100  sub	r4, r0, r4
  448=>x"8861",	-- 1000100001100001  brige	r4, PaperGameQuit
  449=>x"D210",	-- 1101001000010000  sw	r0, r2
  450=>x"0412",	-- 0000010000010010  inc	r2, r2
  451=>x"041B",	-- 0000010000011011  inc	r3, r3
  452=>x"D010",	-- 1101000000010000  lw	r0, r2
  453=>x"D019",	-- 1101000000011001  lw	r1, r3
  454=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  455=>x"D210",	-- 1101001000010000  sw	r0, r2
  456=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  457=>x"1800",	-- 0001100000000000  
  458=>x"D01B",	-- 1101000000011011  lw	r3, r3
  459=>x"BAD8",	-- 1011101011011000  brieq	r3, PaperGameLoop
  460=>x"F7DC",	-- 1111011111011100  bspl	r4, r3, 15
  461=>x"8524",	-- 1000010100100100  brine	r4, PaperGameQuit
  462=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  463=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveUp
  464=>x"F49C",	-- 1111010010011100  bspl	r4, r3, 2
  465=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveDOWN
  466=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  467=>x"81A0",	-- 1000000110100000  brieq	r4, PaperNoMoveLEFT
  468=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  469=>x"173D",	-- 0001011100111101  
  470=>x"D010",	-- 1101000000010000  lw	r0, r2
  471=>x"0600",	-- 0000011000000000  dec	r0, r0
  472=>x"D210",	-- 1101001000010000  sw	r0, r2
  473=>x"F4DC",	-- 1111010011011100  bspl	r4, r3, 3
  474=>x"81A0",	-- 1000000110100000  brieq	r4, PaperNoMoveRIGHT
  475=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  476=>x"173D",	-- 0001011100111101  
  477=>x"D010",	-- 1101000000010000  lw	r0, r2
  478=>x"0400",	-- 0000010000000000  inc	r0, r0
  479=>x"D210",	-- 1101001000010000  sw	r0, r2
  480=>x"A503",	-- 1010010100000011  bri	-, PaperGameRedrawContent
  481=>x"FFFF",	-- 1111111111111111  reset
  482=>x"063F",	-- 0000011000111111  dec	r7, r7
  483=>x"D238",	-- 1101001000111000  sw	r0, r7
  484=>x"063F",	-- 0000011000111111  dec	r7, r7
  485=>x"D239",	-- 1101001000111001  sw	r1, r7
  486=>x"063F",	-- 0000011000111111  dec	r7, r7
  487=>x"D23A",	-- 1101001000111010  sw	r2, r7
  488=>x"063F",	-- 0000011000111111  dec	r7, r7
  489=>x"D23B",	-- 1101001000111011  sw	r3, r7
  490=>x"063F",	-- 0000011000111111  dec	r7, r7
  491=>x"D23C",	-- 1101001000111100  sw	r4, r7
  492=>x"063F",	-- 0000011000111111  dec	r7, r7
  493=>x"D23D",	-- 1101001000111101  sw	r5, r7
  494=>x"063F",	-- 0000011000111111  dec	r7, r7
  495=>x"D23E",	-- 1101001000111110  sw	r6, r7
  496=>x"FFF2",	-- 1111111111110010  liw	r2, paper_tiles
  497=>x"1730",	-- 0001011100110000  
  498=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  499=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  500=>x"C043",	-- 1100000001000011  li	r3, 8
  501=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  502=>x"02BA",	-- 0000001010111010  
  503=>x"D03E",	-- 1101000000111110  lw	r6, r7
  504=>x"043F",	-- 0000010000111111  inc	r7, r7
  505=>x"D03D",	-- 1101000000111101  lw	r5, r7
  506=>x"043F",	-- 0000010000111111  inc	r7, r7
  507=>x"D03C",	-- 1101000000111100  lw	r4, r7
  508=>x"043F",	-- 0000010000111111  inc	r7, r7
  509=>x"D03B",	-- 1101000000111011  lw	r3, r7
  510=>x"043F",	-- 0000010000111111  inc	r7, r7
  511=>x"D03A",	-- 1101000000111010  lw	r2, r7
  512=>x"043F",	-- 0000010000111111  inc	r7, r7
  513=>x"D039",	-- 1101000000111001  lw	r1, r7
  514=>x"043F",	-- 0000010000111111  inc	r7, r7
  515=>x"D038",	-- 1101000000111000  lw	r0, r7
  516=>x"043F",	-- 0000010000111111  inc	r7, r7
  517=>x"0400",	-- 0000010000000000  inc	r0, r0
  518=>x"E383",	-- 1110001110000011  ba	-, r6
  519=>x"C750",	-- 1100011101010000  li	r0, 234
  520=>x"C1C2",	-- 1100000111000010  li	r2, 56
  521=>x"FAC6",	-- 1111101011000110  bail	-, r6, div_16_16
  522=>x"021F",	-- 0000001000011111  
  523=>x"C448",	-- 1100010001001000  li	r0, 137
  524=>x"C472",	-- 1100010001110010  li	r2, 142
  525=>x"FAC6",	-- 1111101011000110  bail	-, r6, mult_16_16
  526=>x"0213",	-- 0000001000010011  
  527=>x"C03A",	-- 1100000000111010  li r2, 7
  528=>x"FAC6",	-- 1111101011000110  bail	-, r6, fact_16
  529=>x"022A",	-- 0000001000101010  
  530=>x"FFFF",	-- 1111111111111111  reset
  531=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  532=>x"2524",	-- 0010010100100100  xor	r4, r4, r4
  533=>x"C085",	-- 1100000010000101  li	r5, 16
  534=>x"0849",	-- 0000100001001001  add	r1, r1, r1
  535=>x"0C00",	-- 0000110000000000  adc	r0, r0, r0
  536=>x"0EDB",	-- 0000111011011011  sbc	r3, r3, r3
  537=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  538=>x"08C9",	-- 0000100011001001  add	r1, r1, r3
  539=>x"0D00",	-- 0000110100000000  adc	r0, r0, r4
  540=>x"062D",	-- 0000011000101101  dec	r5, r5
  541=>x"BE6C",	-- 1011111001101100  brine	r5, mult_16_16.loop
  542=>x"E383",	-- 1110001110000011  ba	-, r6
  543=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  544=>x"C084",	-- 1100000010000100  li	r4, 16
  545=>x"0800",	-- 0000100000000000  add	r0, r0, r0
  546=>x"0C49",	-- 0000110001001001  adc	r1, r1, r1
  547=>x"0A8B",	-- 0000101010001011  sub	r3, r1, r2
  548=>x"80DD",	-- 1000000011011101  brilt	r3, div_16_16.skip
  549=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  550=>x"0400",	-- 0000010000000000  inc	r0, r0
  551=>x"0624",	-- 0000011000100100  dec	r4, r4
  552=>x"BE64",	-- 1011111001100100  brine	r4, div_16_16.loop
  553=>x"E383",	-- 1110001110000011  ba	-, r6
  554=>x"2400",	-- 0010010000000000  xor	r0, r0, r0
  555=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  556=>x"8250",	-- 1000001001010000  brieq	r2, fact_16.end
  557=>x"0409",	-- 0000010000001001  inc	r1, r1
  558=>x"1008",	-- 0001000000001000  mova	r0, r1
  559=>x"FAC6",	-- 1111101011000110  bail	-, r6, mult_16_16
  560=>x"0213",	-- 0000001000010011  
  561=>x"8104",	-- 1000000100000100  brine	r0, fact_16.overflow
  562=>x"0213",	-- 0000001000010011  
  563=>x"0612",	-- 0000011000010010  dec	r2, r2
  564=>x"BE94",	-- 1011111010010100  brine	r2, fact_16.loop
  565=>x"E383",	-- 1110001110000011  ba	-, r6
  566=>x"063F",	-- 0000011000111111  dec	r7, r7
  567=>x"D23E",	-- 1101001000111110  sw	r6, r7
  568=>x"D013",	-- 1101000000010011  lw	r3, r2
  569=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  570=>x"84D8",	-- 1000010011011000  brieq	r3, puts.end
  571=>x"063F",	-- 0000011000111111  dec	r7, r7
  572=>x"D23A",	-- 1101001000111010  sw	r2, r7
  573=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  574=>x"0250",	-- 0000001001010000  
  575=>x"D03A",	-- 1101000000111010  lw	r2, r7
  576=>x"043F",	-- 0000010000111111  inc	r7, r7
  577=>x"D013",	-- 1101000000010011  lw	r3, r2
  578=>x"4E1B",	-- 0100111000011011  shl	r3, r3, 7
  579=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  580=>x"8258",	-- 1000001001011000  brieq	r3, puts.end
  581=>x"063F",	-- 0000011000111111  dec	r7, r7
  582=>x"D23A",	-- 1101001000111010  sw	r2, r7
  583=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  584=>x"0250",	-- 0000001001010000  
  585=>x"D03A",	-- 1101000000111010  lw	r2, r7
  586=>x"043F",	-- 0000010000111111  inc	r7, r7
  587=>x"0412",	-- 0000010000010010  inc	r2, r2
  588=>x"BB03",	-- 1011101100000011  bri	-, puts.loop
  589=>x"D03E",	-- 1101000000111110  lw	r6, r7
  590=>x"043F",	-- 0000010000111111  inc	r7, r7
  591=>x"E383",	-- 1110001110000011  ba	-, r6
  592=>x"063F",	-- 0000011000111111  dec	r7, r7
  593=>x"D23E",	-- 1101001000111110  sw	r6, r7
  594=>x"063F",	-- 0000011000111111  dec	r7, r7
  595=>x"D238",	-- 1101001000111000  sw	r0, r7
  596=>x"063F",	-- 0000011000111111  dec	r7, r7
  597=>x"D239",	-- 1101001000111001  sw	r1, r7
  598=>x"FFF2",	-- 1111111111110010  liw	r2, font_map
  599=>x"12C0",	-- 0001001011000000  
  600=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  601=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  602=>x"C043",	-- 1100000001000011  li	r3, 8
  603=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  604=>x"02BA",	-- 0000001010111010  
  605=>x"D039",	-- 1101000000111001  lw	r1, r7
  606=>x"043F",	-- 0000010000111111  inc	r7, r7
  607=>x"D038",	-- 1101000000111000  lw	r0, r7
  608=>x"043F",	-- 0000010000111111  inc	r7, r7
  609=>x"0400",	-- 0000010000000000  inc	r0, r0
  610=>x"D03E",	-- 1101000000111110  lw	r6, r7
  611=>x"043F",	-- 0000010000111111  inc	r7, r7
  612=>x"E383",	-- 1110001110000011  ba	-, r6
  613=>x"063F",	-- 0000011000111111  dec	r7, r7
  614=>x"D23E",	-- 1101001000111110  sw	r6, r7
  615=>x"FFF4",	-- 1111111111110100  liw	r4, 10000
  616=>x"2710",	-- 0010011100010000  
  617=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  618=>x"0278",	-- 0000001001111000  
  619=>x"FFF4",	-- 1111111111110100  liw	r4, 1000
  620=>x"03E8",	-- 0000001111101000  
  621=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  622=>x"0278",	-- 0000001001111000  
  623=>x"C324",	-- 1100001100100100  li	r4, 100
  624=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  625=>x"0278",	-- 0000001001111000  
  626=>x"C054",	-- 1100000001010100  li	r4, 10
  627=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  628=>x"0278",	-- 0000001001111000  
  629=>x"D03E",	-- 1101000000111110  lw	r6, r7
  630=>x"043F",	-- 0000010000111111  inc	r7, r7
  631=>x"C00C",	-- 1100000000001100  li	r4, 1
  632=>x"C17B",	-- 1100000101111011  li	r3, 0x2F
  633=>x"041B",	-- 0000010000011011  inc	r3, r3
  634=>x"0B12",	-- 0000101100010010  sub	r2, r2, r4
  635=>x"BF91",	-- 1011111110010001  brige	r2, printnum.loop
  636=>x"0912",	-- 0000100100010010  add	r2, r2, r4
  637=>x"063F",	-- 0000011000111111  dec	r7, r7
  638=>x"D23E",	-- 1101001000111110  sw	r6, r7
  639=>x"063F",	-- 0000011000111111  dec	r7, r7
  640=>x"D23A",	-- 1101001000111010  sw	r2, r7
  641=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  642=>x"0250",	-- 0000001001010000  
  643=>x"D03A",	-- 1101000000111010  lw	r2, r7
  644=>x"043F",	-- 0000010000111111  inc	r7, r7
  645=>x"D03E",	-- 1101000000111110  lw	r6, r7
  646=>x"043F",	-- 0000010000111111  inc	r7, r7
  647=>x"E383",	-- 1110001110000011  ba	-, r6
  648=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  649=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  650=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  651=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  652=>x"C0A0",	-- 1100000010100000  li	r0, 20
  653=>x"D011",	-- 1101000000010001  lw	r1, r2
  654=>x"D221",	-- 1101001000100001  sw	r1, r4
  655=>x"0412",	-- 0000010000010010  inc	r2, r2
  656=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  657=>x"061B",	-- 0000011000011011  dec	r3, r3
  658=>x"BEDC",	-- 1011111011011100  brine	r3, put_sprite_16_aligned.loop
  659=>x"E383",	-- 1110001110000011  ba	-, r6
  660=>x"C07D",	-- 1100000001111101  li	r5, 15
  661=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  662=>x"6600",	-- 0110011000000000  shr	r0, r0, 3
  663=>x"BC68",	-- 1011110001101000  brieq	r5, put_sprite_16_aligned
  664=>x"062D",	-- 0000011000101101  dec	r5, r5
  665=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  666=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  667=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  668=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  669=>x"063F",	-- 0000011000111111  dec	r7, r7
  670=>x"D23B",	-- 1101001000111011  sw	r3, r7
  671=>x"D011",	-- 1101000000010001  lw	r1, r2
  672=>x"CFF8",	-- 1100111111111000  li	r0, -1
  673=>x"3D40",	-- 0011110101000000  rsr	r0, r0, r5
  674=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  675=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  676=>x"D023",	-- 1101000000100011  lw	r3, r4
  677=>x"2600",	-- 0010011000000000  not	r0, r0
  678=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  679=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  680=>x"D221",	-- 1101001000100001  sw	r1, r4
  681=>x"0424",	-- 0000010000100100  inc	r4, r4
  682=>x"D011",	-- 1101000000010001  lw	r1, r2
  683=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  684=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  685=>x"D023",	-- 1101000000100011  lw	r3, r4
  686=>x"2600",	-- 0010011000000000  not	r0, r0
  687=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  688=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  689=>x"D221",	-- 1101001000100001  sw	r1, r4
  690=>x"0412",	-- 0000010000010010  inc	r2, r2
  691=>x"C098",	-- 1100000010011000  li	r0, 19
  692=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  693=>x"D03B",	-- 1101000000111011  lw	r3, r7
  694=>x"043F",	-- 0000010000111111  inc	r7, r7
  695=>x"061B",	-- 0000011000011011  dec	r3, r3
  696=>x"B95C",	-- 1011100101011100  brine	r3, put_sprite_16.loop
  697=>x"E383",	-- 1110001110000011  ba	-, r6
  698=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  699=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  700=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  701=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  702=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  703=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  704=>x"C0A5",	-- 1100000010100101  li	r5, 20
  705=>x"8404",	-- 1000010000000100  brine	r0, put_sprite_8_aligned.loop1
  706=>x"D010",	-- 1101000000010000  lw	r0, r2
  707=>x"D021",	-- 1101000000100001  lw	r1, r4
  708=>x"1A41",	-- 0001101001000001  mixhl	r1, r0, r1
  709=>x"D221",	-- 1101001000100001  sw	r1, r4
  710=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  711=>x"061B",	-- 0000011000011011  dec	r3, r3
  712=>x"E398",	-- 1110001110011000  baeq	r3, r6
  713=>x"D021",	-- 1101000000100001  lw	r1, r4
  714=>x"1E41",	-- 0001111001000001  mixll	r1, r0, r1
  715=>x"D221",	-- 1101001000100001  sw	r1, r4
  716=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  717=>x"0412",	-- 0000010000010010  inc	r2, r2
  718=>x"061B",	-- 0000011000011011  dec	r3, r3
  719=>x"E398",	-- 1110001110011000  baeq	r3, r6
  720=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop0
  721=>x"D010",	-- 1101000000010000  lw	r0, r2
  722=>x"D021",	-- 1101000000100001  lw	r1, r4
  723=>x"1809",	-- 0001100000001001  mixhh	r1, r1, r0
  724=>x"D221",	-- 1101001000100001  sw	r1, r4
  725=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  726=>x"061B",	-- 0000011000011011  dec	r3, r3
  727=>x"E398",	-- 1110001110011000  baeq	r3, r6
  728=>x"D021",	-- 1101000000100001  lw	r1, r4
  729=>x"1A09",	-- 0001101000001001  mixhl	r1, r1, r0
  730=>x"D221",	-- 1101001000100001  sw	r1, r4
  731=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  732=>x"0412",	-- 0000010000010010  inc	r2, r2
  733=>x"061B",	-- 0000011000011011  dec	r3, r3
  734=>x"E398",	-- 1110001110011000  baeq	r3, r6
  735=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop1
  736=>x"C03D",	-- 1100000000111101  li	r5, 7
  737=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  738=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  739=>x"B5E8",	-- 1011010111101000  brieq	r5, put_sprite_8_aligned
  740=>x"062D",	-- 0000011000101101  dec	r5, r5
  741=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  742=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  743=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  744=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  745=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  746=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  747=>x"8A04",	-- 1000101000000100  brine	r0, put_sprite_8.loop1
  748=>x"D010",	-- 1101000000010000  lw	r0, r2
  749=>x"063F",	-- 0000011000111111  dec	r7, r7
  750=>x"D23A",	-- 1101001000111010  sw	r2, r7
  751=>x"C802",	-- 1100100000000010  li	r2, 0x100
  752=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  753=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  754=>x"D021",	-- 1101000000100001  lw	r1, r4
  755=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  756=>x"2612",	-- 0010011000010010  not	r2, r2
  757=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  758=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  759=>x"D221",	-- 1101001000100001  sw	r1, r4
  760=>x"C0A1",	-- 1100000010100001  li	r1, 20
  761=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  762=>x"D03A",	-- 1101000000111010  lw	r2, r7
  763=>x"043F",	-- 0000010000111111  inc	r7, r7
  764=>x"061B",	-- 0000011000011011  dec	r3, r3
  765=>x"E398",	-- 1110001110011000  baeq	r3, r6
  766=>x"D010",	-- 1101000000010000  lw	r0, r2
  767=>x"063F",	-- 0000011000111111  dec	r7, r7
  768=>x"D23A",	-- 1101001000111010  sw	r2, r7
  769=>x"1E00",	-- 0001111000000000  mixll	r0, r0, r0
  770=>x"C802",	-- 1100100000000010  li	r2, 0x100
  771=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  772=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  773=>x"D021",	-- 1101000000100001  lw	r1, r4
  774=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  775=>x"2612",	-- 0010011000010010  not	r2, r2
  776=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  777=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  778=>x"D221",	-- 1101001000100001  sw	r1, r4
  779=>x"C0A1",	-- 1100000010100001  li	r1, 20
  780=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  781=>x"D03A",	-- 1101000000111010  lw	r2, r7
  782=>x"043F",	-- 0000010000111111  inc	r7, r7
  783=>x"0412",	-- 0000010000010010  inc	r2, r2
  784=>x"061B",	-- 0000011000011011  dec	r3, r3
  785=>x"E398",	-- 1110001110011000  baeq	r3, r6
  786=>x"B683",	-- 1011011010000011  bri	-, put_sprite_8.loop0
  787=>x"D010",	-- 1101000000010000  lw	r0, r2
  788=>x"063F",	-- 0000011000111111  dec	r7, r7
  789=>x"D23A",	-- 1101001000111010  sw	r2, r7
  790=>x"063F",	-- 0000011000111111  dec	r7, r7
  791=>x"D23B",	-- 1101001000111011  sw	r3, r7
  792=>x"C802",	-- 1100100000000010  li	r2, 0x100
  793=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  794=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  795=>x"2080",	-- 0010000010000000  and	r0, r0, r2
  796=>x"D021",	-- 1101000000100001  lw	r1, r4
  797=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
  798=>x"261B",	-- 0010011000011011  not	r3, r3
  799=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  800=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
  801=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  802=>x"D221",	-- 1101001000100001  sw	r1, r4
  803=>x"0424",	-- 0000010000100100  inc	r4, r4
  804=>x"D021",	-- 1101000000100001  lw	r1, r4
  805=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  806=>x"261B",	-- 0010011000011011  not	r3, r3
  807=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  808=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
  809=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  810=>x"D221",	-- 1101001000100001  sw	r1, r4
  811=>x"C099",	-- 1100000010011001  li	r1, 19
  812=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  813=>x"D03B",	-- 1101000000111011  lw	r3, r7
  814=>x"043F",	-- 0000010000111111  inc	r7, r7
  815=>x"D03A",	-- 1101000000111010  lw	r2, r7
  816=>x"043F",	-- 0000010000111111  inc	r7, r7
  817=>x"061B",	-- 0000011000011011  dec	r3, r3
  818=>x"E398",	-- 1110001110011000  baeq	r3, r6
  819=>x"D010",	-- 1101000000010000  lw	r0, r2
  820=>x"4E00",	-- 0100111000000000  shl	r0, r0, 7
  821=>x"063F",	-- 0000011000111111  dec	r7, r7
  822=>x"D23A",	-- 1101001000111010  sw	r2, r7
  823=>x"063F",	-- 0000011000111111  dec	r7, r7
  824=>x"D23B",	-- 1101001000111011  sw	r3, r7
  825=>x"C802",	-- 1100100000000010  li	r2, 0x100
  826=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  827=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  828=>x"2080",	-- 0010000010000000  and	r0, r0, r2
  829=>x"D021",	-- 1101000000100001  lw	r1, r4
  830=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
  831=>x"261B",	-- 0010011000011011  not	r3, r3
  832=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  833=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
  834=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  835=>x"D221",	-- 1101001000100001  sw	r1, r4
  836=>x"0424",	-- 0000010000100100  inc	r4, r4
  837=>x"D021",	-- 1101000000100001  lw	r1, r4
  838=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  839=>x"261B",	-- 0010011000011011  not	r3, r3
  840=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
  841=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
  842=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  843=>x"D221",	-- 1101001000100001  sw	r1, r4
  844=>x"C099",	-- 1100000010011001  li	r1, 19
  845=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  846=>x"D03B",	-- 1101000000111011  lw	r3, r7
  847=>x"043F",	-- 0000010000111111  inc	r7, r7
  848=>x"D03A",	-- 1101000000111010  lw	r2, r7
  849=>x"043F",	-- 0000010000111111  inc	r7, r7
  850=>x"0412",	-- 0000010000010010  inc	r2, r2
  851=>x"061B",	-- 0000011000011011  dec	r3, r3
  852=>x"E398",	-- 1110001110011000  baeq	r3, r6
  853=>x"AF83",	-- 1010111110000011  bri	-, put_sprite_8.loop1
    others => x"0000"
    );
begin
  process(CLK)
  begin
    if (CLK'event AND CLK='1') then
      D <= m(to_integer(unsigned(AD)));
    end if;
  end process;
end Behavioral;
