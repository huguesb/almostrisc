----------------------------------------------------------------------------------
--
-- File retrieved, on 07/02/2010, from :
-- http://sebastien-viardot.imag.fr/Enseignements/Archi1A2s/sources/ROMPROG.vhd
--
-- Slightly altered to get rid of vendor-specific packages and adjust formatting
-- Now auto-filled by asrom script
--
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROMPROG is
  Port ( AD : in  STD_LOGIC_VECTOR (12 downto 0);
         D : out  STD_LOGIC_VECTOR (15 downto 0);
         CLK : in STD_LOGIC);
end ROMPROG;

architecture Behavioral of ROMPROG is
  constant low_address: natural := 0;
  constant high_address: natural := 8192;
  subtype octet is std_logic_vector( 15 downto 0 );
  type zone_memoire is
    array (natural range low_address to high_address-1) of octet;
  constant m: zone_memoire:= (
    0=>x"FFF7",	-- 1111111111110111  liw	r7, IRQ_mask
    1=>x"2000",	-- 0010000000000000  
    2=>x"F8C0",	-- 1111100011000000  bai	-, os_init
    3=>x"0100",	-- 0000000100000000  
   16=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_ack
   17=>x"2002",	-- 0010000000000010  
   18=>x"D001",	-- 1101000000000001  lw	r1, r0
   19=>x"F54A",	-- 1111010101001010  bspl	r2, r1, 5
   20=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_error
   21=>x"0050",	-- 0000000001010000  
   22=>x"F4CA",	-- 1111010011001010  bspl	r2, r1, 3
   23=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_kbd
   24=>x"0060",	-- 0000000001100000  
   25=>x"F40A",	-- 1111010000001010  bspl	r2, r1, 0
   26=>x"FB16",	-- 1111101100010110  bailne	r2, r6, int_tmr
   27=>x"0040",	-- 0000000001000000  
   28=>x"D201",	-- 1101001000000001  sw	r1, r0
   29=>x"FFFE",	-- 1111111111111110  reti
   64=>x"263F",	-- 0010011000111111  not r7, r7
   65=>x"D7C0",	-- 1101011111000000  out	r7
   66=>x"E383",	-- 1110001110000011  ba	-, r6
   80=>x"25FF",	-- 0010010111111111  xor	r7, r7, r7
   81=>x"D7C0",	-- 1101011111000000  out	r7
   82=>x"E383",	-- 1110001110000011  ba	-, r6
   96=>x"FFF2",	-- 1111111111110010  liw	r2, PS2_rx
   97=>x"2004",	-- 0010000000000100  
   98=>x"D012",	-- 1101000000010010  lw	r2, r2
   99=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map + 8
  100=>x"16C8",	-- 0001011011001000  
  101=>x"D01B",	-- 1101000000011011  lw	r3, r3
  102=>x"1EBF",	-- 0001111010111111  mixll	r7, r7, r2
  103=>x"C784",	-- 1100011110000100  li	r4, 0xF0
  104=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  105=>x"8C60",	-- 1000110001100000  brieq	r4, int_kbd.release
  106=>x"C704",	-- 1100011100000100  li	r4, 0xE0
  107=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  108=>x"8A20",	-- 1000101000100000  brieq	r4, int_kbd.extended
  109=>x"FFF5",	-- 1111111111110101  liw	r5, rand_seed
  110=>x"16C8",	-- 0001011011001000  
  111=>x"D02C",	-- 1101000000101100  lw	r4, r5
  112=>x"24A4",	-- 0010010010100100  xor	r4, r4, r2
  113=>x"D22C",	-- 1101001000101100  sw	r4, r5
  114=>x"FFF5",	-- 1111111111110101  liw	r5, paper_keys - 1
  115=>x"16CF",	-- 0001011011001111  
  116=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  117=>x"80E0",	-- 1000000011100000  brieq	r4, $+3
  118=>x"FFF5",	-- 1111111111110101  liw	r5, paper_keys + 11 - 1
  119=>x"16DA",	-- 0001011011011010  
  120=>x"042D",	-- 0000010000101101  inc	r5, r5
  121=>x"D02C",	-- 1101000000101100  lw	r4, r5
  122=>x"8560",	-- 1000010101100000  brieq	r4, scan_code_mismatch
  123=>x"6E24",	-- 0110111000100100  shr	r4, r4, 7
  124=>x"0B14",	-- 0000101100010100  sub	r4, r2, r4
  125=>x"BEE4",	-- 1011111011100100  brine	r4, scan_code_loop
  126=>x"D02A",	-- 1101000000101010  lw	r2, r5
  127=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  128=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
  129=>x"741B",	-- 0111010000011011  shr	r3, r3, 10
  130=>x"C00D",	-- 1100000000001101  li	r5, 1
  131=>x"0612",	-- 0000011000010010  dec	r2, r2
  132=>x"3AAA",	-- 0011101010101010  rrl	r2, r5, r2
  133=>x"FFF5",	-- 1111111111110101  liw	r5, key_press_map
  134=>x"16C0",	-- 0001011011000000  
  135=>x"08ED",	-- 0000100011101101  add	r5, r5, r3
  136=>x"D02B",	-- 1101000000101011  lw	r3, r5
  137=>x"80E4",	-- 1000000011100100  brine	r4, scan_code_release
  138=>x"229B",	-- 0010001010011011  or	r3, r3, r2
  139=>x"80C3",	-- 1000000011000011  bri	-, scan_code_notify
  140=>x"2612",	-- 0010011000010010  not	r2, r2
  141=>x"209B",	-- 0010000010011011  and	r3, r3, r2
  142=>x"D22B",	-- 1101001000101011  sw	r3, r5
  143=>x"C003",	-- 1100000000000011  li	r3, 0
  144=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  145=>x"16C8",	-- 0001011011001000  
  146=>x"D223",	-- 1101001000100011  sw	r3, r4
  147=>x"E383",	-- 1110001110000011  ba	-, r6
  148=>x"C014",	-- 1100000000010100  li	r4, 2
  149=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  150=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  151=>x"16C8",	-- 0001011011001000  
  152=>x"D223",	-- 1101001000100011  sw	r3, r4
  153=>x"E383",	-- 1110001110000011  ba	-, r6
  154=>x"C00C",	-- 1100000000001100  li	r4, 1
  155=>x"231B",	-- 0010001100011011  or	r3, r3, r4
  156=>x"FFF4",	-- 1111111111110100  liw	r4, key_press_map + 8
  157=>x"16C8",	-- 0001011011001000  
  158=>x"D223",	-- 1101001000100011  sw	r3, r4
  159=>x"E383",	-- 1110001110000011  ba	-, r6
  256=>x"FFF0",	-- 1111111111110000  liw	r0, IRQ_mask
  257=>x"2000",	-- 0010000000000000  
  258=>x"C0C9",	-- 1100000011001001  li	r1, 0x19
  259=>x"D201",	-- 1101001000000001  sw	r1, r0
  260=>x"0400",	-- 0000010000000000  inc	r0, r0
  261=>x"CFF9",	-- 1100111111111001  li	r1, -1
  262=>x"D201",	-- 1101001000000001  sw	r1, r0
  263=>x"C03A",	-- 1100000000111010  li	r2, 7
  264=>x"0880",	-- 0000100010000000  add	r0, r0, r2
  265=>x"C0EA",	-- 1100000011101010  li	r2, 0x1D
  266=>x"D202",	-- 1101001000000010  sw	r2, r0
  267=>x"0400",	-- 0000010000000000  inc	r0, r0
  268=>x"C07A",	-- 1100000001111010  li	r2, 15
  269=>x"D202",	-- 1101001000000010  sw	r2, r0
  270=>x"0400",	-- 0000010000000000  inc	r0, r0
  271=>x"C0DA",	-- 1100000011011010  li	r2, 0x1B
  272=>x"D202",	-- 1101001000000010  sw	r2, r0
  273=>x"0400",	-- 0000010000000000  inc	r0, r0
  274=>x"FFF2",	-- 1111111111110010  liw	r2, 817
  275=>x"0331",	-- 0000001100110001  
  276=>x"D202",	-- 1101001000000010  sw	r2, r0
  277=>x"FFF0",	-- 1111111111110000  liw	r0, key_press_map
  278=>x"16C0",	-- 0001011011000000  
  279=>x"C001",	-- 1100000000000001  li	r1, 0
  280=>x"C042",	-- 1100000001000010  li	r2, 8
  281=>x"D201",	-- 1101001000000001  sw	r1, r0
  282=>x"0400",	-- 0000010000000000  inc	r0, r0
  283=>x"0612",	-- 0000011000010010  dec	r2, r2
  284=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  285=>x"8083",	-- 1000000010000011  bri	-, PaperGameStart
  286=>x"8003",	-- 1000000000000011  bri	-, PaperMenuLoop
  287=>x"FFF0",	-- 1111111111110000  liw	r0, paper_score
  288=>x"16C9",	-- 0001011011001001  
  289=>x"C001",	-- 1100000000000001  li	r1, 0
  290=>x"D201",	-- 1101001000000001  sw	r1, r0
  291=>x"FFF0",	-- 1111111111110000  liw	r0, paper_dir
  292=>x"179C",	-- 0001011110011100  
  293=>x"C001",	-- 1100000000000001  li	r1, 0
  294=>x"D201",	-- 1101001000000001  sw	r1, r0
  295=>x"0400",	-- 0000010000000000  inc	r0, r0
  296=>x"FFF1",	-- 1111111111110001  liw	r1, 152 * 8
  297=>x"04C0",	-- 0000010011000000  
  298=>x"D201",	-- 1101001000000001  sw	r1, r0
  299=>x"0400",	-- 0000010000000000  inc	r0, r0
  300=>x"C001",	-- 1100000000000001  li	r1, 0
  301=>x"D201",	-- 1101001000000001  sw	r1, r0
  302=>x"0400",	-- 0000010000000000  inc	r0, r0
  303=>x"FFF1",	-- 1111111111110001  liw	r1, 128 * 8
  304=>x"0400",	-- 0000010000000000  
  305=>x"D201",	-- 1101001000000001  sw	r1, r0
  306=>x"0400",	-- 0000010000000000  inc	r0, r0
  307=>x"C001",	-- 1100000000000001  li	r1, 0
  308=>x"D201",	-- 1101001000000001  sw	r1, r0
  309=>x"0400",	-- 0000010000000000  inc	r0, r0
  310=>x"C069",	-- 1100000001101001  li	r1, 13
  311=>x"D201",	-- 1101001000000001  sw	r1, r0
  312=>x"0400",	-- 0000010000000000  inc	r0, r0
  313=>x"C011",	-- 1100000000010001  li	r1, 2
  314=>x"D201",	-- 1101001000000001  sw	r1, r0
  315=>x"0400",	-- 0000010000000000  inc	r0, r0
  316=>x"FFF0",	-- 1111111111110000  liw	r0, paper_tilemap
  317=>x"17B0",	-- 0001011110110000  
  318=>x"C001",	-- 1100000000000001  li	r1, 0
  319=>x"C0C2",	-- 1100000011000010  li	r2, 6*4
  320=>x"D201",	-- 1101001000000001  sw	r1, r0
  321=>x"0400",	-- 0000010000000000  inc	r0, r0
  322=>x"0612",	-- 0000011000010010  dec	r2, r2
  323=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  324=>x"C000",	-- 1100000000000000  li	r0, 0
  325=>x"CFF9",	-- 1100111111111001  li	r1, -1
  326=>x"C0A2",	-- 1100000010100010  li	r2, 20
  327=>x"D201",	-- 1101001000000001  sw	r1, r0
  328=>x"0400",	-- 0000010000000000  inc	r0, r0
  329=>x"0612",	-- 0000011000010010  dec	r2, r2
  330=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  331=>x"C001",	-- 1100000000000001  li	r1, 0
  332=>x"FFF2",	-- 1111111111110010  liw	r2, 18*20
  333=>x"0168",	-- 0000000101101000  
  334=>x"D201",	-- 1101001000000001  sw	r1, r0
  335=>x"0400",	-- 0000010000000000  inc	r0, r0
  336=>x"0612",	-- 0000011000010010  dec	r2, r2
  337=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  338=>x"CFF9",	-- 1100111111111001  li	r1, -1
  339=>x"C0A2",	-- 1100000010100010  li	r2, 20
  340=>x"D201",	-- 1101001000000001  sw	r1, r0
  341=>x"0400",	-- 0000010000000000  inc	r0, r0
  342=>x"0612",	-- 0000011000010010  dec	r2, r2
  343=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  344=>x"C020",	-- 1100000000100000  li	r0, 4
  345=>x"C029",	-- 1100000000101001  li	r1, 5
  346=>x"FFF2",	-- 1111111111110010  liw	r2, paper_title
  347=>x"17A4",	-- 0001011110100100  
  348=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  349=>x"02BF",	-- 0000001010111111  
  350=>x"C090",	-- 1100000010010000  li	r0, 18
  351=>x"C029",	-- 1100000000101001  li	r1, 5
  352=>x"FFF2",	-- 1111111111110010  liw	r2, paper_score
  353=>x"16C9",	-- 0001011011001001  
  354=>x"D012",	-- 1101000000010010  lw	r2, r2
  355=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum
  356=>x"02EE",	-- 0000001011101110  
  357=>x"C778",	-- 1100011101111000  li	r0, 239
  358=>x"C009",	-- 1100000000001001  li	r1, 1
  359=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud
  360=>x"1780",	-- 0001011110000000  
  361=>x"C043",	-- 1100000001000011  li	r3, 8
  362=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  363=>x"03C7",	-- 0000001111000111  
  364=>x"C0F8",	-- 1100000011111000  li	r0, 31
  365=>x"C009",	-- 1100000000001001  li	r1, 1
  366=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  367=>x"17A0",	-- 0001011110100000  
  368=>x"D012",	-- 1101000000010010  lw	r2, r2
  369=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum
  370=>x"02EE",	-- 0000001011101110  
  371=>x"C120",	-- 1100000100100000  li	r0, 36
  372=>x"C009",	-- 1100000000001001  li	r1, 1
  373=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  374=>x"17AA",	-- 0001011110101010  
  375=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  376=>x"02BF",	-- 0000001010111111  
  377=>x"C778",	-- 1100011101111000  li	r0, 239
  378=>x"C051",	-- 1100000001010001  li	r1, 10
  379=>x"FFF2",	-- 1111111111110010  liw	r2, paper_hud + 8
  380=>x"1788",	-- 0001011110001000  
  381=>x"C043",	-- 1100000001000011  li	r3, 8
  382=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8
  383=>x"03C7",	-- 0000001111000111  
  384=>x"C0F8",	-- 1100000011111000  li	r0, 31
  385=>x"C051",	-- 1100000001010001  li	r1, 10
  386=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed + 1
  387=>x"17A1",	-- 0001011110100001  
  388=>x"D012",	-- 1101000000010010  lw	r2, r2
  389=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum
  390=>x"02EE",	-- 0000001011101110  
  391=>x"C120",	-- 1100000100100000  li	r0, 36
  392=>x"C051",	-- 1100000001010001  li	r1, 10
  393=>x"FFF2",	-- 1111111111110010  liw	r2, paper_unit
  394=>x"17AA",	-- 0001011110101010  
  395=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  396=>x"02BF",	-- 0000001010111111  
  397=>x"FFF0",	-- 1111111111110000  liw	r0, 20*20
  398=>x"0190",	-- 0000000110010000  
  399=>x"C001",	-- 1100000000000001  li	r1, 0
  400=>x"FFF2",	-- 1111111111110010  liw	r2, 220*20
  401=>x"1130",	-- 0001000100110000  
  402=>x"D201",	-- 1101001000000001  sw	r1, r0
  403=>x"0400",	-- 0000010000000000  inc	r0, r0
  404=>x"0612",	-- 0000011000010010  dec	r2, r2
  405=>x"BF54",	-- 1011111101010100  brine	r2, $-3
  406=>x"FFF5",	-- 1111111111110101  liw	r5, paper_tilemap
  407=>x"17B0",	-- 0001011110110000  
  408=>x"D02C",	-- 1101000000101100  lw	r4, r5
  409=>x"042D",	-- 0000010000101101  inc	r5, r5
  410=>x"8960",	-- 1000100101100000  brieq	r4, PaperGameTileSkip
  411=>x"063F",	-- 0000011000111111  dec	r7, r7
  412=>x"D23D",	-- 1101001000111101  sw	r5, r7
  413=>x"FFF3",	-- 1111111111110011  liw	r3, paper_tilemap
  414=>x"17B0",	-- 0001011110110000  
  415=>x"0AEB",	-- 0000101011101011  sub	r3, r5, r3
  416=>x"6E20",	-- 0110111000100000  shr	r0, r4, 7
  417=>x"6219",	-- 0110001000011001  shr	r1, r3, 1
  418=>x"4809",	-- 0100100000001001  shl	r1, r1, 4
  419=>x"C19A",	-- 1100000110011010  li	r2, 51
  420=>x"0889",	-- 0000100010001001  add	r1, r1, r2
  421=>x"FFF2",	-- 1111111111110010  liw	r2, paper_pos + 1
  422=>x"179E",	-- 0001011110011110  
  423=>x"D012",	-- 1101000000010010  lw	r2, r2
  424=>x"6412",	-- 0110010000010010  shr	r2, r2, 2
  425=>x"C0FB",	-- 1100000011111011  li	r3, 31
  426=>x"20D2",	-- 0010000011010010  and	r2, r2, r3
  427=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  428=>x"4E24",	-- 0100111000100100  shl	r4, r4, 7
  429=>x"6E24",	-- 0110111000100100  shr	r4, r4, 7
  430=>x"C00B",	-- 1100000000001011  li	r3, 1
  431=>x"FB06",	-- 1111101100000110  bailne	r0, r6, put_tile
  432=>x"028F",	-- 0000001010001111  
  433=>x"81E0",	-- 1000000111100000  brieq	r4, PaperGameSegmentSkip
  435=>x"C013",	-- 1100000000010011  li	r3, 2
  436=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_tile
  437=>x"028F",	-- 0000001010001111  
  438=>x"0624",	-- 0000011000100100  dec	r4, r4
  439=>x"BF64",	-- 1011111101100100  brine	r4, PaperGameSegmentLoop
  440=>x"C003",	-- 1100000000000011  li	r3, 0
  441=>x"C144",	-- 1100000101000100  li	r4, 40
  442=>x"0B04",	-- 0000101100000100  sub	r4, r0, r4
  443=>x"FB66",	-- 1111101101100110  baillt	r4, r6, put_tile
  444=>x"028F",	-- 0000001010001111  
  445=>x"D03D",	-- 1101000000111101  lw	r5, r7
  446=>x"043F",	-- 0000010000111111  inc	r7, r7
  447=>x"FFF4",	-- 1111111111110100  liw r4, paper_tilemap + 24
  448=>x"17C8",	-- 0001011111001000  
  449=>x"0B2C",	-- 0000101100101100  sub	r4, r5, r4
  450=>x"B5A5",	-- 1011010110100101  brilt	r4, PaperGameTileLoop
  451=>x"FFF3",	-- 1111111111110011  liw	r3, paper_speed
  452=>x"17A0",	-- 0001011110100000  
  453=>x"D01B",	-- 1101000000011011  lw	r3, r3
  454=>x"CF04",	-- 1100111100000100  li	r4, 0x1E0
  455=>x"211C",	-- 0010000100011100  and	r4, r3, r4
  456=>x"FFF3",	-- 1111111111110011  liw	r3, paper_pos
  457=>x"179D",	-- 0001011110011101  
  458=>x"D018",	-- 1101000000011000  lw	r0, r3
  459=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  460=>x"FFF2",	-- 1111111111110010  liw	r2, paper_sprites
  461=>x"1720",	-- 0001011100100000  
  462=>x"0912",	-- 0000100100010010  add	r2, r2, r4
  463=>x"C161",	-- 1100000101100001  li	r1, 44
  464=>x"C083",	-- 1100000010000011  li	r3, 16
  465=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_16_masked
  466=>x"035F",	-- 0000001101011111  
  467=>x"90AC",	-- 1001000010101100  brine	r5, PaperGameFail
  469=>x"C028",	-- 1100000000101000  li	r0, 5
  470=>x"C001",	-- 1100000000000001  li	r1, 0
  471=>x"8043",	-- 1000000001000011  bri	-, $+1
  472=>x"0609",	-- 0000011000001001  dec	r1, r1
  473=>x"BF8C",	-- 1011111110001100  brine	r1, $-2
  474=>x"0600",	-- 0000011000000000  dec	r0, r0
  475=>x"BEC4",	-- 1011111011000100  brine	r0, $-5
  476=>x"FFF2",	-- 1111111111110010  liw	r2, paper_pos
  477=>x"179D",	-- 0001011110011101  
  478=>x"FFF3",	-- 1111111111110011  liw	r3, paper_speed
  479=>x"17A0",	-- 0001011110100000  
  480=>x"D010",	-- 1101000000010000  lw	r0, r2
  481=>x"D019",	-- 1101000000011001  lw	r1, r3
  482=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  483=>x"8C85",	-- 1000110010000101  brilt	r0, PaperGameFail
  484=>x"FFF4",	-- 1111111111110100  liw	r4, 304*8
  485=>x"0980",	-- 0000100110000000  
  486=>x"0B04",	-- 0000101100000100  sub	r4, r0, r4
  487=>x"8BA1",	-- 1000101110100001  brige	r4, PaperGameFail
  488=>x"D210",	-- 1101001000010000  sw	r0, r2
  489=>x"0412",	-- 0000010000010010  inc	r2, r2
  490=>x"041B",	-- 0000010000011011  inc	r3, r3
  491=>x"D010",	-- 1101000000010000  lw	r0, r2
  492=>x"D019",	-- 1101000000011001  lw	r1, r3
  493=>x"C7FC",	-- 1100011111111100  li	r4, 0xFF
  494=>x"6009",	-- 0110000000001001  shr	r1, r1, 0
  495=>x"0840",	-- 0000100001000000  add	r0, r0, r1
  496=>x"2101",	-- 0010000100000001  and	r1, r0, r4
  497=>x"D211",	-- 1101001000010001  sw	r1, r2
  498=>x"2624",	-- 0010011000100100  not	r4, r4
  499=>x"2100",	-- 0010000100000000  and	r0, r0, r4
  500=>x"FB06",	-- 1111101100000110  bailne	r0, r6, PaperMapScroll
  501=>x"0237",	-- 0000001000110111  
  502=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  503=>x"16C0",	-- 0001011011000000  
  504=>x"D01B",	-- 1101000000011011  lw	r3, r3
  505=>x"F818",	-- 1111100000011000  baieq	r3, PaperGameRedraw
  506=>x"0144",	-- 0000000101000100  
  507=>x"F55C",	-- 1111010101011100  bspl	r4, r3, 5
  508=>x"8AA4",	-- 1000101010100100  brine	r4, PaperGameQuit
  509=>x"F51C",	-- 1111010100011100  bspl	r4, r3, 4
  510=>x"8A64",	-- 1000101001100100  brine	r4, PaperGamePause
  511=>x"F41C",	-- 1111010000011100  bspl	r4, r3, 0
  512=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveUp
  513=>x"F49C",	-- 1111010010011100  bspl	r4, r3, 2
  514=>x"8060",	-- 1000000001100000  brieq	r4, PaperNoMoveDOWN
  515=>x"F45C",	-- 1111010001011100  bspl	r4, r3, 1
  516=>x"81E0",	-- 1000000111100000  brieq	r4, PaperNoMoveLEFT
  517=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  518=>x"17A0",	-- 0001011110100000  
  519=>x"D010",	-- 1101000000010000  lw	r0, r2
  520=>x"C02C",	-- 1100000000101100  li	r4, 5
  521=>x"0B00",	-- 0000101100000000  sub	r0, r0, r4
  522=>x"D210",	-- 1101001000010000  sw	r0, r2
  523=>x"F4DC",	-- 1111010011011100  bspl	r4, r3, 3
  524=>x"81E0",	-- 1000000111100000  brieq	r4, PaperNoMoveRIGHT
  525=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed
  526=>x"17A0",	-- 0001011110100000  
  527=>x"D010",	-- 1101000000010000  lw	r0, r2
  528=>x"C02C",	-- 1100000000101100  li	r4, 5
  529=>x"0900",	-- 0000100100000000  add	r0, r0, r4
  530=>x"D210",	-- 1101001000010000  sw	r0, r2
  531=>x"F8C0",	-- 1111100011000000  bai	-, PaperGameRedraw
  532=>x"0144",	-- 0000000101000100  
  533=>x"C000",	-- 1100000000000000  li	r0, 0
  534=>x"FFF2",	-- 1111111111110010  liw	r2, 240*20
  535=>x"12C0",	-- 0001001011000000  
  536=>x"D001",	-- 1101000000000001  lw	r1, r0
  537=>x"2609",	-- 0010011000001001  not	r1, r1
  538=>x"D201",	-- 1101001000000001  sw	r1, r0
  539=>x"0400",	-- 0000010000000000  inc	r0, r0
  540=>x"0612",	-- 0000011000010010  dec	r2, r2
  541=>x"BED4",	-- 1011111011010100  brine	r2, $-5
  542=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  543=>x"16C0",	-- 0001011011000000  
  544=>x"D01A",	-- 1101000000011010  lw	r2, r3
  545=>x"BFD4",	-- 1011111111010100  brine	r2, $-1
  546=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  547=>x"16C0",	-- 0001011011000000  
  548=>x"D01A",	-- 1101000000011010  lw	r2, r3
  549=>x"BFD0",	-- 1011111111010000  brieq	r2, $-1
  550=>x"FFFF",	-- 1111111111111111  reset
  551=>x"C080",	-- 1100000010000000  li	r0, 16
  552=>x"C0C1",	-- 1100000011000001  li	r1, 24
  553=>x"FFF2",	-- 1111111111110010  liw	r2, paper_pause
  554=>x"17C8",	-- 0001011111001000  
  555=>x"FAC6",	-- 1111101011000110  bail	-, r6, puts
  556=>x"02BF",	-- 0000001010111111  
  557=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  558=>x"16C0",	-- 0001011011000000  
  559=>x"D01A",	-- 1101000000011010  lw	r2, r3
  560=>x"BFD4",	-- 1011111111010100  brine	r2, $-1
  561=>x"FFF3",	-- 1111111111110011  liw	r3, key_press_map
  562=>x"16C0",	-- 0001011011000000  
  563=>x"D01A",	-- 1101000000011010  lw	r2, r3
  564=>x"BFD0",	-- 1011111111010000  brieq	r2, $-1
  565=>x"F8C0",	-- 1111100011000000  bai	-, PaperGameRedraw
  566=>x"0144",	-- 0000000101000100  
  567=>x"FFF0",	-- 1111111111110000  liw	r0, paper_tilemap
  568=>x"17B0",	-- 0001011110110000  
  569=>x"C021",	-- 1100000000100001  li	r1, 4
  570=>x"0841",	-- 0000100001000001  add	r1, r0, r1
  571=>x"C0A2",	-- 1100000010100010  li	r2, 5*4
  572=>x"D00B",	-- 1101000000001011  lw	r3, r1
  573=>x"D203",	-- 1101001000000011  sw	r3, r0
  574=>x"0400",	-- 0000010000000000  inc	r0, r0
  575=>x"0409",	-- 0000010000001001  inc	r1, r1
  576=>x"0612",	-- 0000011000010010  dec	r2, r2
  577=>x"BED4",	-- 1011111011010100  brine	r2, PaperGameScrollLoop
  578=>x"063F",	-- 0000011000111111  dec	r7, r7
  579=>x"D23E",	-- 1101001000111110  sw	r6, r7
  580=>x"FAC6",	-- 1111101011000110  bail	-, r6, rand16
  581=>x"027D",	-- 0000001001111101  
  582=>x"C02A",	-- 1100000000101010  li	r2, 0x05
  583=>x"208B",	-- 0010000010001011  and	r3, r1, r2
  584=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  585=>x"208C",	-- 0010000010001100  and	r4, r1, r2
  586=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  587=>x"1F19",	-- 0001111100011001  mixll	r1, r3, r4
  588=>x"D201",	-- 1101001000000001  sw	r1, r0
  589=>x"0400",	-- 0000010000000000  inc	r0, r0
  590=>x"C03A",	-- 1100000000111010  li	r2, 0x07
  591=>x"091C",	-- 0000100100011100  add r4, r3, r4
  592=>x"208B",	-- 0010000010001011  and	r3, r1, r2
  593=>x"091C",	-- 0000100100011100  add r4, r3, r4
  594=>x"C01B",	-- 1100000000011011  li	r3, 3
  595=>x"08E4",	-- 0000100011100100  add	r4, r4, r3
  596=>x"6209",	-- 0110001000001001  shr	r1, r1, 1
  597=>x"208B",	-- 0010000010001011  and	r3, r1, r2
  598=>x"091B",	-- 0000100100011011  add r3, r3, r4
  599=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  600=>x"208C",	-- 0010000010001100  and	r4, r1, r2
  601=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  602=>x"1F19",	-- 0001111100011001  mixll	r1, r3, r4
  603=>x"D201",	-- 1101001000000001  sw	r1, r0
  604=>x"0400",	-- 0000010000000000  inc	r0, r0
  605=>x"C02A",	-- 1100000000101010  li	r2, 0x05
  606=>x"091C",	-- 0000100100011100  add r4, r3, r4
  607=>x"208B",	-- 0010000010001011  and	r3, r1, r2
  608=>x"091C",	-- 0000100100011100  add r4, r3, r4
  609=>x"C01B",	-- 1100000000011011  li	r3, 3
  610=>x"08E4",	-- 0000100011100100  add	r4, r4, r3
  611=>x"6209",	-- 0110001000001001  shr	r1, r1, 1
  612=>x"208B",	-- 0010000010001011  and	r3, r1, r2
  613=>x"091B",	-- 0000100100011011  add r3, r3, r4
  614=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  615=>x"208C",	-- 0010000010001100  and	r4, r1, r2
  616=>x"6409",	-- 0110010000001001  shr	r1, r1, 2
  617=>x"1F19",	-- 0001111100011001  mixll	r1, r3, r4
  618=>x"D201",	-- 1101001000000001  sw	r1, r0
  619=>x"0400",	-- 0000010000000000  inc	r0, r0
  620=>x"FFF2",	-- 1111111111110010  liw	r2, paper_speed + 1
  621=>x"17A1",	-- 0001011110100001  
  622=>x"D011",	-- 1101000000010001  lw	r1, r2
  623=>x"0409",	-- 0000010000001001  inc	r1, r1
  624=>x"D211",	-- 1101001000010001  sw	r1, r2
  625=>x"FFF2",	-- 1111111111110010  liw	r2, paper_score
  626=>x"16C9",	-- 0001011011001001  
  627=>x"D011",	-- 1101000000010001  lw	r1, r2
  628=>x"0409",	-- 0000010000001001  inc	r1, r1
  629=>x"D211",	-- 1101001000010001  sw	r1, r2
  630=>x"D03E",	-- 1101000000111110  lw	r6, r7
  631=>x"043F",	-- 0000010000111111  inc	r7, r7
  632=>x"E383",	-- 1110001110000011  ba	-, r6
  633=>x"FFF2",	-- 1111111111110010  liw	r2, rand_seed
  634=>x"16C8",	-- 0001011011001000  
  635=>x"D210",	-- 1101001000010000  sw	r0, r2
  636=>x"E383",	-- 1110001110000011  ba	-, r6
  637=>x"FFF2",	-- 1111111111110010  liw	r2, rand_seed
  638=>x"16C8",	-- 0001011011001000  
  639=>x"D013",	-- 1101000000010011  lw	r3, r2
  640=>x"C7EC",	-- 1100011111101100  li	r4, 253
  641=>x"1F19",	-- 0001111100011001  mixll	r1, r3, r4
  642=>x"18E4",	-- 0001100011100100  mixhh	r4, r4, r3
  643=>x"C002",	-- 1100000000000010  li	r2, 0
  644=>x"0AC9",	-- 0000101011001001  sub	r1, r1, r3
  645=>x"0EA4",	-- 0000111010100100  sbc	r4, r4, r2
  646=>x"0EC9",	-- 0000111011001001  sbc	r1, r1, r3
  647=>x"0EA4",	-- 0000111010100100  sbc	r4, r4, r2
  648=>x"1B13",	-- 0001101100010011  mixhl	r3, r2, r4
  649=>x"0EC9",	-- 0000111011001001  sbc	r1, r1, r3
  650=>x"0C89",	-- 0000110010001001  adc	r1, r1, r2
  651=>x"FFF2",	-- 1111111111110010  liw	r2, rand_seed
  652=>x"16C8",	-- 0001011011001000  
  653=>x"D211",	-- 1101001000010001  sw	r1, r2
  654=>x"E383",	-- 1110001110000011  ba	-, r6
  655=>x"063F",	-- 0000011000111111  dec	r7, r7
  656=>x"D238",	-- 1101001000111000  sw	r0, r7
  657=>x"063F",	-- 0000011000111111  dec	r7, r7
  658=>x"D239",	-- 1101001000111001  sw	r1, r7
  659=>x"063F",	-- 0000011000111111  dec	r7, r7
  660=>x"D23A",	-- 1101001000111010  sw	r2, r7
  661=>x"063F",	-- 0000011000111111  dec	r7, r7
  662=>x"D23B",	-- 1101001000111011  sw	r3, r7
  663=>x"063F",	-- 0000011000111111  dec	r7, r7
  664=>x"D23C",	-- 1101001000111100  sw	r4, r7
  665=>x"063F",	-- 0000011000111111  dec	r7, r7
  666=>x"D23D",	-- 1101001000111101  sw	r5, r7
  667=>x"063F",	-- 0000011000111111  dec	r7, r7
  668=>x"D23E",	-- 1101001000111110  sw	r6, r7
  669=>x"FFF2",	-- 1111111111110010  liw	r2, paper_tiles
  670=>x"1790",	-- 0001011110010000  
  671=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  672=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  673=>x"C043",	-- 1100000001000011  li	r3, 8
  674=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  675=>x"03A1",	-- 0000001110100001  
  676=>x"D03E",	-- 1101000000111110  lw	r6, r7
  677=>x"043F",	-- 0000010000111111  inc	r7, r7
  678=>x"D03D",	-- 1101000000111101  lw	r5, r7
  679=>x"043F",	-- 0000010000111111  inc	r7, r7
  680=>x"D03C",	-- 1101000000111100  lw	r4, r7
  681=>x"043F",	-- 0000010000111111  inc	r7, r7
  682=>x"D03B",	-- 1101000000111011  lw	r3, r7
  683=>x"043F",	-- 0000010000111111  inc	r7, r7
  684=>x"D03A",	-- 1101000000111010  lw	r2, r7
  685=>x"043F",	-- 0000010000111111  inc	r7, r7
  686=>x"D039",	-- 1101000000111001  lw	r1, r7
  687=>x"043F",	-- 0000010000111111  inc	r7, r7
  688=>x"D038",	-- 1101000000111000  lw	r0, r7
  689=>x"043F",	-- 0000010000111111  inc	r7, r7
  690=>x"0400",	-- 0000010000000000  inc	r0, r0
  691=>x"E383",	-- 1110001110000011  ba	-, r6
  692=>x"2449",	-- 0010010001001001  xor	r1, r1, r1
  693=>x"C084",	-- 1100000010000100  li	r4, 16
  694=>x"0800",	-- 0000100000000000  add	r0, r0, r0
  695=>x"0C49",	-- 0000110001001001  adc	r1, r1, r1
  696=>x"0A8B",	-- 0000101010001011  sub	r3, r1, r2
  697=>x"80DD",	-- 1000000011011101  brilt	r3, div_16_16.skip
  698=>x"0A89",	-- 0000101010001001  sub	r1, r1, r2
  699=>x"0400",	-- 0000010000000000  inc	r0, r0
  700=>x"0624",	-- 0000011000100100  dec	r4, r4
  701=>x"BE64",	-- 1011111001100100  brine	r4, div_16_16.loop
  702=>x"E383",	-- 1110001110000011  ba	-, r6
  703=>x"063F",	-- 0000011000111111  dec	r7, r7
  704=>x"D23E",	-- 1101001000111110  sw	r6, r7
  705=>x"D013",	-- 1101000000010011  lw	r3, r2
  706=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  707=>x"84D8",	-- 1000010011011000  brieq	r3, puts.end
  708=>x"063F",	-- 0000011000111111  dec	r7, r7
  709=>x"D23A",	-- 1101001000111010  sw	r2, r7
  710=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  711=>x"02D9",	-- 0000001011011001  
  712=>x"D03A",	-- 1101000000111010  lw	r2, r7
  713=>x"043F",	-- 0000010000111111  inc	r7, r7
  714=>x"D013",	-- 1101000000010011  lw	r3, r2
  715=>x"4E1B",	-- 0100111000011011  shl	r3, r3, 7
  716=>x"6E1B",	-- 0110111000011011  shr	r3, r3, 7
  717=>x"8258",	-- 1000001001011000  brieq	r3, puts.end
  718=>x"063F",	-- 0000011000111111  dec	r7, r7
  719=>x"D23A",	-- 1101001000111010  sw	r2, r7
  720=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  721=>x"02D9",	-- 0000001011011001  
  722=>x"D03A",	-- 1101000000111010  lw	r2, r7
  723=>x"043F",	-- 0000010000111111  inc	r7, r7
  724=>x"0412",	-- 0000010000010010  inc	r2, r2
  725=>x"BB03",	-- 1011101100000011  bri	-, puts.loop
  726=>x"D03E",	-- 1101000000111110  lw	r6, r7
  727=>x"043F",	-- 0000010000111111  inc	r7, r7
  728=>x"E383",	-- 1110001110000011  ba	-, r6
  729=>x"063F",	-- 0000011000111111  dec	r7, r7
  730=>x"D23E",	-- 1101001000111110  sw	r6, r7
  731=>x"063F",	-- 0000011000111111  dec	r7, r7
  732=>x"D238",	-- 1101001000111000  sw	r0, r7
  733=>x"063F",	-- 0000011000111111  dec	r7, r7
  734=>x"D239",	-- 1101001000111001  sw	r1, r7
  735=>x"FFF2",	-- 1111111111110010  liw	r2, font_map
  736=>x"12C0",	-- 0001001011000000  
  737=>x"421B",	-- 0100001000011011  shl	r3, r3, 1
  738=>x"08D2",	-- 0000100011010010  add	r2, r2, r3
  739=>x"C043",	-- 1100000001000011  li	r3, 8
  740=>x"FAC6",	-- 1111101011000110  bail	-, r6, put_sprite_8_aligned
  741=>x"03A1",	-- 0000001110100001  
  742=>x"D039",	-- 1101000000111001  lw	r1, r7
  743=>x"043F",	-- 0000010000111111  inc	r7, r7
  744=>x"D038",	-- 1101000000111000  lw	r0, r7
  745=>x"043F",	-- 0000010000111111  inc	r7, r7
  746=>x"0400",	-- 0000010000000000  inc	r0, r0
  747=>x"D03E",	-- 1101000000111110  lw	r6, r7
  748=>x"043F",	-- 0000010000111111  inc	r7, r7
  749=>x"E383",	-- 1110001110000011  ba	-, r6
  750=>x"063F",	-- 0000011000111111  dec	r7, r7
  751=>x"D23E",	-- 1101001000111110  sw	r6, r7
  752=>x"FFF4",	-- 1111111111110100  liw	r4, 10000
  753=>x"2710",	-- 0010011100010000  
  754=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  755=>x"0301",	-- 0000001100000001  
  756=>x"FFF4",	-- 1111111111110100  liw	r4, 1000
  757=>x"03E8",	-- 0000001111101000  
  758=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  759=>x"0301",	-- 0000001100000001  
  760=>x"C324",	-- 1100001100100100  li	r4, 100
  761=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  762=>x"0301",	-- 0000001100000001  
  763=>x"C054",	-- 1100000001010100  li	r4, 10
  764=>x"FAC6",	-- 1111101011000110  bail	-, r6, printnum.sub
  765=>x"0301",	-- 0000001100000001  
  766=>x"D03E",	-- 1101000000111110  lw	r6, r7
  767=>x"043F",	-- 0000010000111111  inc	r7, r7
  768=>x"C00C",	-- 1100000000001100  li	r4, 1
  769=>x"C17B",	-- 1100000101111011  li	r3, 0x2F
  770=>x"041B",	-- 0000010000011011  inc	r3, r3
  771=>x"0B12",	-- 0000101100010010  sub	r2, r2, r4
  772=>x"BF91",	-- 1011111110010001  brige	r2, printnum.loop
  773=>x"0912",	-- 0000100100010010  add	r2, r2, r4
  774=>x"063F",	-- 0000011000111111  dec	r7, r7
  775=>x"D23E",	-- 1101001000111110  sw	r6, r7
  776=>x"063F",	-- 0000011000111111  dec	r7, r7
  777=>x"D23A",	-- 1101001000111010  sw	r2, r7
  778=>x"FAC6",	-- 1111101011000110  bail	-, r6, putchar
  779=>x"02D9",	-- 0000001011011001  
  780=>x"D03A",	-- 1101000000111010  lw	r2, r7
  781=>x"043F",	-- 0000010000111111  inc	r7, r7
  782=>x"D03E",	-- 1101000000111110  lw	r6, r7
  783=>x"043F",	-- 0000010000111111  inc	r7, r7
  784=>x"E383",	-- 1110001110000011  ba	-, r6
  785=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  786=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  787=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  788=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  789=>x"C0A0",	-- 1100000010100000  li	r0, 20
  790=>x"0412",	-- 0000010000010010  inc	r2, r2
  791=>x"D011",	-- 1101000000010001  lw	r1, r2
  792=>x"E421",	-- 1110010000100001  exw	r1, r4
  793=>x"0412",	-- 0000010000010010  inc	r2, r2
  794=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  795=>x"061B",	-- 0000011000011011  dec	r3, r3
  796=>x"BE9C",	-- 1011111010011100  brine	r3, put_sprite_16_aligned.loop
  797=>x"C005",	-- 1100000000000101  li	r5, 0
  798=>x"E383",	-- 1110001110000011  ba	-, r6
  799=>x"C07D",	-- 1100000001111101  li	r5, 15
  800=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  801=>x"6600",	-- 0110011000000000  shr	r0, r0, 3
  802=>x"BBE8",	-- 1011101111101000  brieq	r5, put_sprite_16_aligned
  803=>x"062D",	-- 0000011000101101  dec	r5, r5
  804=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  805=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  806=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  807=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  808=>x"063F",	-- 0000011000111111  dec	r7, r7
  809=>x"D23B",	-- 1101001000111011  sw	r3, r7
  810=>x"0412",	-- 0000010000010010  inc	r2, r2
  811=>x"D011",	-- 1101000000010001  lw	r1, r2
  812=>x"CFF8",	-- 1100111111111000  li	r0, -1
  813=>x"3D40",	-- 0011110101000000  rsr	r0, r0, r5
  814=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  815=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  816=>x"D023",	-- 1101000000100011  lw	r3, r4
  817=>x"2600",	-- 0010011000000000  not	r0, r0
  818=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  819=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  820=>x"E421",	-- 1110010000100001  exw	r1, r4
  821=>x"0424",	-- 0000010000100100  inc	r4, r4
  822=>x"D011",	-- 1101000000010001  lw	r1, r2
  823=>x"3949",	-- 0011100101001001  rrr	r1, r1, r5
  824=>x"2009",	-- 0010000000001001  and	r1, r1, r0
  825=>x"D023",	-- 1101000000100011  lw	r3, r4
  826=>x"2600",	-- 0010011000000000  not	r0, r0
  827=>x"201B",	-- 0010000000011011  and	r3, r3, r0
  828=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
  829=>x"E421",	-- 1110010000100001  exw	r1, r4
  830=>x"0412",	-- 0000010000010010  inc	r2, r2
  831=>x"C098",	-- 1100000010011000  li	r0, 19
  832=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  833=>x"D03B",	-- 1101000000111011  lw	r3, r7
  834=>x"043F",	-- 0000010000111111  inc	r7, r7
  835=>x"061B",	-- 0000011000011011  dec	r3, r3
  836=>x"B91C",	-- 1011100100011100  brine	r3, put_sprite_16.loop
  837=>x"C005",	-- 1100000000000101  li	r5, 0
  838=>x"E383",	-- 1110001110000011  ba	-, r6
  839=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  840=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  841=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  842=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  843=>x"C005",	-- 1100000000000101  li	r5, 0
  844=>x"D020",	-- 1101000000100000  lw	r0, r4
  845=>x"D011",	-- 1101000000010001  lw	r1, r2
  846=>x"0412",	-- 0000010000010010  inc	r2, r2
  847=>x"2040",	-- 0010000001000000  and	r0, r0, r1
  848=>x"D011",	-- 1101000000010001  lw	r1, r2
  849=>x"2240",	-- 0010001001000000  or	r0, r0, r1
  850=>x"E420",	-- 1110010000100000  exw	r0, r4
  851=>x"0612",	-- 0000011000010010  dec	r2, r2
  852=>x"D011",	-- 1101000000010001  lw	r1, r2
  853=>x"2609",	-- 0010011000001001  not	r1, r1
  854=>x"0412",	-- 0000010000010010  inc	r2, r2
  855=>x"2040",	-- 0010000001000000  and	r0, r0, r1
  856=>x"222D",	-- 0010001000101101  or	r5, r5, r0
  857=>x"0412",	-- 0000010000010010  inc	r2, r2
  858=>x"C0A0",	-- 1100000010100000  li	r0, 20
  859=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  860=>x"061B",	-- 0000011000011011  dec	r3, r3
  861=>x"AE5C",	-- 1010111001011100  brine	r3, put_sprite_16_aligned.loop
  862=>x"E383",	-- 1110001110000011  ba	-, r6
  863=>x"C07D",	-- 1100000001111101  li	r5, 15
  864=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  865=>x"6600",	-- 0110011000000000  shr	r0, r0, 3
  866=>x"B968",	-- 1011100101101000  brieq	r5, put_sprite_16_masked_aligned
  867=>x"062D",	-- 0000011000101101  dec	r5, r5
  868=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  869=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  870=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  871=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  872=>x"063F",	-- 0000011000111111  dec	r7, r7
  873=>x"D23E",	-- 1101001000111110  sw	r6, r7
  874=>x"102E",	-- 0001000000101110  mova	r6, r5
  875=>x"C005",	-- 1100000000000101  li	r5, 0
  876=>x"063F",	-- 0000011000111111  dec	r7, r7
  877=>x"D23B",	-- 1101001000111011  sw	r3, r7
  878=>x"063F",	-- 0000011000111111  dec	r7, r7
  879=>x"D23D",	-- 1101001000111101  sw	r5, r7
  880=>x"D010",	-- 1101000000010000  lw	r0, r2
  881=>x"3980",	-- 0011100110000000  rrr	r0, r0, r6
  882=>x"0412",	-- 0000010000010010  inc	r2, r2
  883=>x"D011",	-- 1101000000010001  lw	r1, r2
  884=>x"3989",	-- 0011100110001001  rrr	r1, r1, r6
  885=>x"CFFD",	-- 1100111111111101  li	r5, -1
  886=>x"3DAD",	-- 0011110110101101  rsr	r5, r5, r6
  887=>x"2149",	-- 0010000101001001  and	r1, r1, r5
  888=>x"D023",	-- 1101000000100011  lw	r3, r4
  889=>x"262D",	-- 0010011000101101  not	r5, r5
  890=>x"222D",	-- 0010001000101101  or	r5, r5, r0
  891=>x"215B",	-- 0010000101011011  and	r3, r3, r5
  892=>x"225B",	-- 0010001001011011  or	r3, r3, r1
  893=>x"E423",	-- 1110010000100011  exw	r3, r4
  894=>x"262D",	-- 0010011000101101  not	r5, r5
  895=>x"215B",	-- 0010000101011011  and	r3, r3, r5
  896=>x"D03D",	-- 1101000000111101  lw	r5, r7
  897=>x"043F",	-- 0000010000111111  inc	r7, r7
  898=>x"22ED",	-- 0010001011101101  or	r5, r5, r3
  899=>x"0424",	-- 0000010000100100  inc	r4, r4
  900=>x"063F",	-- 0000011000111111  dec	r7, r7
  901=>x"D23D",	-- 1101001000111101  sw	r5, r7
  902=>x"D011",	-- 1101000000010001  lw	r1, r2
  903=>x"3989",	-- 0011100110001001  rrr	r1, r1, r6
  904=>x"CFFD",	-- 1100111111111101  li	r5, -1
  905=>x"3DAD",	-- 0011110110101101  rsr	r5, r5, r6
  906=>x"262D",	-- 0010011000101101  not	r5, r5
  907=>x"2149",	-- 0010000101001001  and	r1, r1, r5
  908=>x"D023",	-- 1101000000100011  lw	r3, r4
  909=>x"262D",	-- 0010011000101101  not	r5, r5
  910=>x"222D",	-- 0010001000101101  or	r5, r5, r0
  911=>x"215B",	-- 0010000101011011  and	r3, r3, r5
  912=>x"225B",	-- 0010001001011011  or	r3, r3, r1
  913=>x"E423",	-- 1110010000100011  exw	r3, r4
  914=>x"262D",	-- 0010011000101101  not	r5, r5
  915=>x"215B",	-- 0010000101011011  and	r3, r3, r5
  916=>x"D03D",	-- 1101000000111101  lw	r5, r7
  917=>x"043F",	-- 0000010000111111  inc	r7, r7
  918=>x"22ED",	-- 0010001011101101  or	r5, r5, r3
  919=>x"0412",	-- 0000010000010010  inc	r2, r2
  920=>x"C098",	-- 1100000010011000  li	r0, 19
  921=>x"0824",	-- 0000100000100100  add	r4, r4, r0
  922=>x"D03B",	-- 1101000000111011  lw	r3, r7
  923=>x"043F",	-- 0000010000111111  inc	r7, r7
  924=>x"061B",	-- 0000011000011011  dec	r3, r3
  925=>x"B3DC",	-- 1011001111011100  brine	r3, put_sprite_16_masked.loop
  926=>x"D03E",	-- 1101000000111110  lw	r6, r7
  927=>x"043F",	-- 0000010000111111  inc	r7, r7
  928=>x"E383",	-- 1110001110000011  ba	-, r6
  929=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  930=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  931=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  932=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  933=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  934=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  935=>x"C0A5",	-- 1100000010100101  li	r5, 20
  936=>x"8404",	-- 1000010000000100  brine	r0, put_sprite_8_aligned.loop1
  937=>x"D010",	-- 1101000000010000  lw	r0, r2
  938=>x"D021",	-- 1101000000100001  lw	r1, r4
  939=>x"1A41",	-- 0001101001000001  mixhl	r1, r0, r1
  940=>x"D221",	-- 1101001000100001  sw	r1, r4
  941=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  942=>x"061B",	-- 0000011000011011  dec	r3, r3
  943=>x"E398",	-- 1110001110011000  baeq	r3, r6
  944=>x"D021",	-- 1101000000100001  lw	r1, r4
  945=>x"1E41",	-- 0001111001000001  mixll	r1, r0, r1
  946=>x"D221",	-- 1101001000100001  sw	r1, r4
  947=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  948=>x"0412",	-- 0000010000010010  inc	r2, r2
  949=>x"061B",	-- 0000011000011011  dec	r3, r3
  950=>x"E398",	-- 1110001110011000  baeq	r3, r6
  951=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop0
  952=>x"D010",	-- 1101000000010000  lw	r0, r2
  953=>x"D021",	-- 1101000000100001  lw	r1, r4
  954=>x"1809",	-- 0001100000001001  mixhh	r1, r1, r0
  955=>x"D221",	-- 1101001000100001  sw	r1, r4
  956=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  957=>x"061B",	-- 0000011000011011  dec	r3, r3
  958=>x"E398",	-- 1110001110011000  baeq	r3, r6
  959=>x"D021",	-- 1101000000100001  lw	r1, r4
  960=>x"1A09",	-- 0001101000001001  mixhl	r1, r1, r0
  961=>x"D221",	-- 1101001000100001  sw	r1, r4
  962=>x"0964",	-- 0000100101100100  add	r4, r4, r5
  963=>x"0412",	-- 0000010000010010  inc	r2, r2
  964=>x"061B",	-- 0000011000011011  dec	r3, r3
  965=>x"E398",	-- 1110001110011000  baeq	r3, r6
  966=>x"BC83",	-- 1011110010000011  bri	-, put_sprite_8_aligned.loop1
  967=>x"C03D",	-- 1100000000111101  li	r5, 7
  968=>x"2145",	-- 0010000101000101  and	r5, r0, r5
  969=>x"6400",	-- 0110010000000000  shr	r0, r0, 2
  970=>x"B5E8",	-- 1011010111101000  brieq	r5, put_sprite_8_aligned
  971=>x"062D",	-- 0000011000101101  dec	r5, r5
  972=>x"460C",	-- 0100011000001100  shl r4, r1, 3
  973=>x"4209",	-- 0100001000001001  shl	r1, r1, 1
  974=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  975=>x"6001",	-- 0110000000000001  shr	r1, r0, 0
  976=>x"0E00",	-- 0000111000000000  sbc	r0, r0, r0
  977=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  978=>x"8A04",	-- 1000101000000100  brine	r0, put_sprite_8.loop1
  979=>x"D010",	-- 1101000000010000  lw	r0, r2
  980=>x"063F",	-- 0000011000111111  dec	r7, r7
  981=>x"D23A",	-- 1101001000111010  sw	r2, r7
  982=>x"C802",	-- 1100100000000010  li	r2, 0x100
  983=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
  984=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
  985=>x"D021",	-- 1101000000100001  lw	r1, r4
  986=>x"2010",	-- 0010000000010000  and	r0, r2, r0
  987=>x"2612",	-- 0010011000010010  not	r2, r2
  988=>x"2089",	-- 0010000010001001  and	r1, r1, r2
  989=>x"2209",	-- 0010001000001001  or	r1, r1, r0
  990=>x"D221",	-- 1101001000100001  sw	r1, r4
  991=>x"C0A1",	-- 1100000010100001  li	r1, 20
  992=>x"0864",	-- 0000100001100100  add	r4, r4, r1
  993=>x"D03A",	-- 1101000000111010  lw	r2, r7
  994=>x"043F",	-- 0000010000111111  inc	r7, r7
  995=>x"061B",	-- 0000011000011011  dec	r3, r3
  996=>x"E398",	-- 1110001110011000  baeq	r3, r6
  997=>x"D010",	-- 1101000000010000  lw	r0, r2
  998=>x"063F",	-- 0000011000111111  dec	r7, r7
  999=>x"D23A",	-- 1101001000111010  sw	r2, r7
 1000=>x"1E00",	-- 0001111000000000  mixll	r0, r0, r0
 1001=>x"C802",	-- 1100100000000010  li	r2, 0x100
 1002=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
 1003=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
 1004=>x"D021",	-- 1101000000100001  lw	r1, r4
 1005=>x"2010",	-- 0010000000010000  and	r0, r2, r0
 1006=>x"2612",	-- 0010011000010010  not	r2, r2
 1007=>x"2089",	-- 0010000010001001  and	r1, r1, r2
 1008=>x"2209",	-- 0010001000001001  or	r1, r1, r0
 1009=>x"D221",	-- 1101001000100001  sw	r1, r4
 1010=>x"C0A1",	-- 1100000010100001  li	r1, 20
 1011=>x"0864",	-- 0000100001100100  add	r4, r4, r1
 1012=>x"D03A",	-- 1101000000111010  lw	r2, r7
 1013=>x"043F",	-- 0000010000111111  inc	r7, r7
 1014=>x"0412",	-- 0000010000010010  inc	r2, r2
 1015=>x"061B",	-- 0000011000011011  dec	r3, r3
 1016=>x"E398",	-- 1110001110011000  baeq	r3, r6
 1017=>x"B683",	-- 1011011010000011  bri	-, put_sprite_8.loop0
 1018=>x"D010",	-- 1101000000010000  lw	r0, r2
 1019=>x"063F",	-- 0000011000111111  dec	r7, r7
 1020=>x"D23A",	-- 1101001000111010  sw	r2, r7
 1021=>x"063F",	-- 0000011000111111  dec	r7, r7
 1022=>x"D23B",	-- 1101001000111011  sw	r3, r7
 1023=>x"C802",	-- 1100100000000010  li	r2, 0x100
 1024=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
 1025=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
 1026=>x"2080",	-- 0010000010000000  and	r0, r0, r2
 1027=>x"D021",	-- 1101000000100001  lw	r1, r4
 1028=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
 1029=>x"261B",	-- 0010011000011011  not	r3, r3
 1030=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
 1031=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
 1032=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
 1033=>x"D221",	-- 1101001000100001  sw	r1, r4
 1034=>x"0424",	-- 0000010000100100  inc	r4, r4
 1035=>x"D021",	-- 1101000000100001  lw	r1, r4
 1036=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
 1037=>x"261B",	-- 0010011000011011  not	r3, r3
 1038=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
 1039=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
 1040=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
 1041=>x"D221",	-- 1101001000100001  sw	r1, r4
 1042=>x"C099",	-- 1100000010011001  li	r1, 19
 1043=>x"0864",	-- 0000100001100100  add	r4, r4, r1
 1044=>x"D03B",	-- 1101000000111011  lw	r3, r7
 1045=>x"043F",	-- 0000010000111111  inc	r7, r7
 1046=>x"D03A",	-- 1101000000111010  lw	r2, r7
 1047=>x"043F",	-- 0000010000111111  inc	r7, r7
 1048=>x"061B",	-- 0000011000011011  dec	r3, r3
 1049=>x"E398",	-- 1110001110011000  baeq	r3, r6
 1050=>x"D010",	-- 1101000000010000  lw	r0, r2
 1051=>x"4E00",	-- 0100111000000000  shl	r0, r0, 7
 1052=>x"063F",	-- 0000011000111111  dec	r7, r7
 1053=>x"D23A",	-- 1101001000111010  sw	r2, r7
 1054=>x"063F",	-- 0000011000111111  dec	r7, r7
 1055=>x"D23B",	-- 1101001000111011  sw	r3, r7
 1056=>x"C802",	-- 1100100000000010  li	r2, 0x100
 1057=>x"3952",	-- 0011100101010010  rrr	r2, r2, r5
 1058=>x"3940",	-- 0011100101000000  rrr	r0, r0, r5
 1059=>x"2080",	-- 0010000010000000  and	r0, r0, r2
 1060=>x"D021",	-- 1101000000100001  lw	r1, r4
 1061=>x"6E13",	-- 0110111000010011  shr	r3, r2, 7
 1062=>x"261B",	-- 0010011000011011  not	r3, r3
 1063=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
 1064=>x"6E03",	-- 0110111000000011  shr	r3, r0, 7
 1065=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
 1066=>x"D221",	-- 1101001000100001  sw	r1, r4
 1067=>x"0424",	-- 0000010000100100  inc	r4, r4
 1068=>x"D021",	-- 1101000000100001  lw	r1, r4
 1069=>x"4E13",	-- 0100111000010011  shl	r3, r2, 7
 1070=>x"261B",	-- 0010011000011011  not	r3, r3
 1071=>x"20C9",	-- 0010000011001001  and	r1, r1, r3
 1072=>x"4E03",	-- 0100111000000011  shl	r3, r0, 7
 1073=>x"22C9",	-- 0010001011001001  or	r1, r1, r3
 1074=>x"D221",	-- 1101001000100001  sw	r1, r4
 1075=>x"C099",	-- 1100000010011001  li	r1, 19
 1076=>x"0864",	-- 0000100001100100  add	r4, r4, r1
 1077=>x"D03B",	-- 1101000000111011  lw	r3, r7
 1078=>x"043F",	-- 0000010000111111  inc	r7, r7
 1079=>x"D03A",	-- 1101000000111010  lw	r2, r7
 1080=>x"043F",	-- 0000010000111111  inc	r7, r7
 1081=>x"0412",	-- 0000010000010010  inc	r2, r2
 1082=>x"061B",	-- 0000011000011011  dec	r3, r3
 1083=>x"E398",	-- 1110001110011000  baeq	r3, r6
 1084=>x"AF83",	-- 1010111110000011  bri	-, put_sprite_8.loop1
    others => x"0000"
    );
begin
  process(CLK)
  begin
    if (CLK'event AND CLK='1') then
      D <= m(to_integer(unsigned(AD)));
    end if;
  end process;
end Behavioral;
